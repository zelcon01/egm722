netcdf S5P_OFFL_L2__CH4____20240407T123946_20240407T142117_33598_03_020600_20240409T045638 {

// global attributes:
		:Conventions = "CF-1.7" ;
		:institution = "KNMI/SRON" ;
		:source = "Sentinel 5 precursor, TROPOMI, space-borne remote sensing, L2" ;
		:history = "2024-04-09 12:47:23 f_s5pops tropnll2dp /mnt/data1/storage_offl_l2/cache_offl_l2/WORKING-613063452/JobOrder.613063423.xml" ;
		:summary = "TROPOMI/S5P Methane 1-Orbit L2 Swath 5.5x7.0km" ;
		:tracking_id = "868827cb-901d-48e7-b9fa-a6d807e5e0c9" ;
		:id = "S5P_OFFL_L2__CH4____20240407T123946_20240407T142117_33598_03_020600_20240409T045638" ;
		:time_reference = "2024-04-07T00:00:00Z" ;
		:time_reference_days_since_1950 = 27125 ;
		:time_reference_julian_day = 2460407.5 ;
		:time_reference_seconds_since_1970 = 1712448000LL ;
		:time_coverage_start = "2024-04-07T13:01:21Z" ;
		:time_coverage_end = "2024-04-07T13:53:37Z" ;
		:time_coverage_duration = "PT3136.488S" ;
		:time_coverage_resolution = "PT0.840S" ;
		:orbit = 33598 ;
		:references = "https://sentinels.copernicus.eu/web/sentinel/technical-guides/sentinel-5p/products-algorithms; http://www.tropomi.eu/data-products/methane" ;
		:processor_version = "2.6.0" ;
		:keywords_vocabulary = "AGU index terms, http://publications.agu.org/author-resource-center/index-terms/" ;
		:keywords = "0300 Atmospheric Composition and Structure; 0365 Troposphere, Composition and Chemistry; 0400 Biogeosciences; 0428 Carbon Cycling; 1600 Global Change" ;
		:standard_name_vocabulary = "NetCDF Climate and Forecast Metadata Conventions Standard Name Table (v29, 08 July 2015), http://cfconventions.org/standard-names.html" ;
		:naming_authority = "nl.knmi" ;
		:cdm_data_type = "Swath" ;
		:date_created = "2024-04-09T05:04:45Z" ;
		:creator_name = "The Sentinel 5 Precursor TROPOMI Level 2 products are developed with funding from the European Space Agency (ESA), the Netherlands Space Office (NSO), the Belgian Science Policy Office, the German Aerospace Center (DLR) and the Bayerisches Staatsministerium für Wirtschaft und Medien, Energie und Technologie (StMWi)." ;
		:creator_url = "https://sentinels.copernicus.eu/web/sentinel/missions/sentinel-5p" ;
		:creator_email = "EOSupport@Copernicus.esa.int" ;
		:project = "Sentinel 5 precursor/TROPOMI" ;
		:geospatial_lat_min = -89.94071f ;
		:geospatial_lat_max = 89.94537f ;
		:geospatial_lon_min = -179.9215f ;
		:geospatial_lon_max = 179.9852f ;
		:license = "No conditions apply" ;
		:platform = "S5P" ;
		:sensor = "TROPOMI" ;
		:spatial_resolution = "5.5x7.0 km2" ;
		:cpp_compiler_version = "g++ (GCC) 4.8.5 20150623 (Red Hat 4.8.5-44)" ;
		:cpp_compiler_flags = "-g -O2 -fPIC -std=c++11 -W -Wall -Wno-ignored-qualifiers -Wno-write-strings -Wno-unused-variable -Wno-unused-parameter -DTROPNLL2DP" ;
		:f90_compiler_version = "GNU Fortran (GCC) 4.8.5 20150623 (Red Hat 4.8.5-44)" ;
		:f90_compiler_flags = "-gdwarf-3 -O2 -fPIC -cpp -ffpe-trap=invalid -fno-range-check -frecursive -fimplicit-none -ffree-line-length-none -DTROPNLL2DP -Wuninitialized -Wtabs" ;
		:build_date = "2023-09-28T07:04:00Z" ;
		:revision_control_identifier = "d084fd110d84" ;
		:geolocation_grid_from_band = 7 ;
		:identifier_product_doi = "10.5270/S5P-3lcdqiv" ;
		:identifier_product_doi_authority = "http://dx.doi.org/" ;
		:algorithm_version = "1.6.0" ;
		:title = "TROPOMI/S5P Methane 1-Orbit L2 Swath 5.5x7.0km" ;
		:product_version = "1.6.0" ;
		:processing_status = "Nominal" ;
		:Status_MET_2D = "Nominal" ;
		:Status_CTM_CO = "Nominal" ;
		:Status_CTMCH4 = "Nominal" ;
		:Status_NPP_VIIRS = "Nominal" ;
		:Status_Internal_Cloud_Mask = "Nominal" ;

group: PRODUCT {
  dimensions:
  	scanline = 3735 ;
  	ground_pixel = 215 ;
  	corner = 4 ;
  	time = 1 ;
  	layer = 12 ;
  	level = 13 ;
  variables:
  	int scanline(scanline) ;
  		scanline:units = "1" ;
  		scanline:axis = "Y" ;
  		scanline:long_name = "along-track dimension index" ;
  		scanline:comment = "This coordinate variable defines the indices along track; index starts at 0" ;
  		scanline:_FillValue = -2147483647 ;
  	int ground_pixel(ground_pixel) ;
  		ground_pixel:units = "1" ;
  		ground_pixel:axis = "X" ;
  		ground_pixel:long_name = "across-track dimension index" ;
  		ground_pixel:comment = "This coordinate variable defines the indices across track, from west to east; index starts at 0" ;
  		ground_pixel:_FillValue = -2147483647 ;
  	int time(time) ;
  		time:units = "seconds since 2010-01-01 00:00:00" ;
  		time:standard_name = "time" ;
  		time:axis = "T" ;
  		time:long_name = "reference time for the measurements" ;
  		time:comment = "The time in this variable corresponds to the time in the time_reference global attribute" ;
  		time:_FillValue = -2147483647 ;
  	int corner(corner) ;
  		corner:units = "1" ;
  		corner:long_name = "pixel corner index" ;
  		corner:comment = "This coordinate variable defines the indices for the pixel corners; index starts at 0 (counter-clockwise, starting from south-western corner of the pixel in ascending part of the orbit)" ;
  		corner:_FillValue = -2147483647 ;
  	int layer(layer) ;
  		layer:axis = "Z" ;
  		layer:positive = "down" ;
  		layer:_FillValue = -2147483647 ;
  	int level(level) ;
  		level:axis = "Z" ;
  		level:positive = "down" ;
  		level:_FillValue = -2147483647 ;
  	int delta_time(time, scanline) ;
  		delta_time:long_name = "offset of start time of measurement relative to time_reference" ;
  		delta_time:units = "milliseconds since 2024-04-07 00:00:00" ;
  		delta_time:_FillValue = -2147483647 ;
  	string time_utc(time, scanline) ;
  		time_utc:long_name = "Time of observation as ISO 8601 date-time string" ;
  		string time_utc:_FillValue = "" ;
  	ubyte qa_value(time, scanline, ground_pixel) ;
  		qa_value:units = "1" ;
  		qa_value:scale_factor = 0.01f ;
  		qa_value:add_offset = 0.f ;
  		qa_value:valid_min = 0UB ;
  		qa_value:valid_max = 100UB ;
  		qa_value:long_name = "data quality value" ;
  		qa_value:comment = "A continuous quality descriptor, varying between 0 (no data) and 1 (full quality data). Recommend to ignore data with qa_value < 0.5" ;
  		qa_value:coordinates = "longitude latitude" ;
  		qa_value:_FillValue = 255UB ;
  	float latitude(time, scanline, ground_pixel) ;
  		latitude:long_name = "pixel center latitude" ;
  		latitude:units = "degrees_north" ;
  		latitude:standard_name = "latitude" ;
  		latitude:valid_min = -90.f ;
  		latitude:valid_max = 90.f ;
  		latitude:bounds = "/PRODUCT/SUPPORT_DATA/GEOLOCATIONS/latitude_bounds" ;
  		latitude:_FillValue = 9.96921e+36f ;
  	float longitude(time, scanline, ground_pixel) ;
  		longitude:long_name = "pixel center longitude" ;
  		longitude:units = "degrees_east" ;
  		longitude:standard_name = "longitude" ;
  		longitude:valid_min = -180.f ;
  		longitude:valid_max = 180.f ;
  		longitude:bounds = "/PRODUCT/SUPPORT_DATA/GEOLOCATIONS/longitude_bounds" ;
  		longitude:_FillValue = 9.96921e+36f ;
  	float methane_mixing_ratio(time, scanline, ground_pixel) ;
  		methane_mixing_ratio:units = "1e-9" ;
  		methane_mixing_ratio:standard_name = "dry_atmosphere_mole_fraction_of_methane" ;
  		methane_mixing_ratio:long_name = "column averaged dry air mixing ratio of methane" ;
  		methane_mixing_ratio:coordinates = "longitude latitude" ;
  		methane_mixing_ratio:ancillary_variables = "methane_mixing_ratio_precision column_averaging_kernel chi_square degreess_of_freedom" ;
  		methane_mixing_ratio:_FillValue = 9.96921e+36f ;
  	float methane_mixing_ratio_precision(time, scanline, ground_pixel) ;
  		methane_mixing_ratio_precision:units = "1e-9" ;
  		methane_mixing_ratio_precision:standard_name = "dry_atmosphere_mole_fraction_of_methane standard_error" ;
  		methane_mixing_ratio_precision:long_name = "precision of the column averaged dry air mixing ratio of methane" ;
  		methane_mixing_ratio_precision:coordinates = "longitude latitude" ;
  		methane_mixing_ratio_precision:_FillValue = 9.96921e+36f ;
  	float methane_mixing_ratio_bias_corrected(time, scanline, ground_pixel) ;
  		methane_mixing_ratio_bias_corrected:units = "1e-9" ;
  		methane_mixing_ratio_bias_corrected:standard_name = "dry_atmosphere_mole_fraction_of_methane" ;
  		methane_mixing_ratio_bias_corrected:long_name = "corrected column-averaged dry-air mole fraction of methane" ;
  		methane_mixing_ratio_bias_corrected:coordinates = "longitude latitude" ;
  		methane_mixing_ratio_bias_corrected:ancillary_variables = "methane_mixing_ratio_precision column_averaging_kernel chi_square degrees_of_freedom" ;
  		methane_mixing_ratio_bias_corrected:comment = "This value will be filled with data after the commissioning phase, this is known to be empty for now" ;
  		methane_mixing_ratio_bias_corrected:_FillValue = 9.96921e+36f ;

  group: SUPPORT_DATA {

    group: GEOLOCATIONS {
      variables:
      	float satellite_latitude(time, scanline) ;
      		satellite_latitude:long_name = "sub satellite latitude" ;
      		satellite_latitude:units = "degrees_north" ;
      		satellite_latitude:comment = "Latitude of the geodetic sub satellite point on the WGS84 reference ellipsoid" ;
      		satellite_latitude:valid_min = -90.f ;
      		satellite_latitude:valid_max = 90.f ;
      		satellite_latitude:_FillValue = 9.96921e+36f ;
      	float satellite_longitude(time, scanline) ;
      		satellite_longitude:long_name = "satellite_longitude" ;
      		satellite_longitude:units = "degrees_east" ;
      		satellite_longitude:comment = "Longitude of the geodetic sub satellite point on the WGS84 reference ellipsoid" ;
      		satellite_longitude:valid_min = -180.f ;
      		satellite_longitude:valid_max = 180.f ;
      		satellite_longitude:_FillValue = 9.96921e+36f ;
      	float satellite_altitude(time, scanline) ;
      		satellite_altitude:long_name = "satellite altitude" ;
      		satellite_altitude:units = "m" ;
      		satellite_altitude:comment = "The altitude of the satellite with respect to the geodetic sub satellite point on the WGS84 reference ellipsoid" ;
      		satellite_altitude:valid_min = 700000.f ;
      		satellite_altitude:valid_max = 900000.f ;
      		satellite_altitude:_FillValue = 9.96921e+36f ;
      	float satellite_orbit_phase(time, scanline) ;
      		satellite_orbit_phase:long_name = "fractional satellite orbit phase" ;
      		satellite_orbit_phase:units = "1" ;
      		satellite_orbit_phase:comment = "Relative offset [0.0, ..., 1.0] of the measurement in the orbit" ;
      		satellite_orbit_phase:valid_min = -0.02f ;
      		satellite_orbit_phase:valid_max = 1.02f ;
      		satellite_orbit_phase:_FillValue = 9.96921e+36f ;
      	float solar_zenith_angle(time, scanline, ground_pixel) ;
      		solar_zenith_angle:long_name = "solar zenith angle" ;
      		solar_zenith_angle:standard_name = "solar_zenith_angle" ;
      		solar_zenith_angle:units = "degree" ;
      		solar_zenith_angle:valid_min = 0.f ;
      		solar_zenith_angle:valid_max = 180.f ;
      		solar_zenith_angle:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		solar_zenith_angle:comment = "Solar zenith angle at the ground pixel location on the reference ellipsoid. Angle is measured away from the vertical" ;
      		solar_zenith_angle:_FillValue = 9.96921e+36f ;
      	float solar_azimuth_angle(time, scanline, ground_pixel) ;
      		solar_azimuth_angle:long_name = "solar azimuth angle" ;
      		solar_azimuth_angle:standard_name = "solar_azimuth_angle" ;
      		solar_azimuth_angle:units = "degree" ;
      		solar_azimuth_angle:valid_min = -180.f ;
      		solar_azimuth_angle:valid_max = 180.f ;
      		solar_azimuth_angle:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		solar_azimuth_angle:comment = "Solar azimuth angle at the ground pixel location on the reference ellipsoid. Angle is measured clockwise from the North (East = 90, South = +/-180, West = -90)" ;
      		solar_azimuth_angle:_FillValue = 9.96921e+36f ;
      	float viewing_zenith_angle(time, scanline, ground_pixel) ;
      		viewing_zenith_angle:long_name = "viewing zenith angle" ;
      		viewing_zenith_angle:standard_name = "viewing_zenith_angle" ;
      		viewing_zenith_angle:units = "degree" ;
      		viewing_zenith_angle:valid_min = 0.f ;
      		viewing_zenith_angle:valid_max = 180.f ;
      		viewing_zenith_angle:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		viewing_zenith_angle:comment = "Zenith angle of the satellite at the ground pixel location on the reference ellipsoid. Angle is measured away from the vertical" ;
      		viewing_zenith_angle:_FillValue = 9.96921e+36f ;
      	float viewing_azimuth_angle(time, scanline, ground_pixel) ;
      		viewing_azimuth_angle:long_name = "viewing azimuth angle" ;
      		viewing_azimuth_angle:standard_name = "viewing_azimuth_angle" ;
      		viewing_azimuth_angle:units = "degree" ;
      		viewing_azimuth_angle:valid_min = -180.f ;
      		viewing_azimuth_angle:valid_max = 180.f ;
      		viewing_azimuth_angle:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		viewing_azimuth_angle:comment = "Satellite azimuth angle at the ground pixel location on the reference ellipsoid. Angle is measured clockwise from the North (East = 90, South = +/-180, West = -90)" ;
      		viewing_azimuth_angle:_FillValue = 9.96921e+36f ;
      	float latitude_bounds(time, scanline, ground_pixel, corner) ;
      		latitude_bounds:_FillValue = 9.96921e+36f ;
      	float longitude_bounds(time, scanline, ground_pixel, corner) ;
      		longitude_bounds:_FillValue = 9.96921e+36f ;
      	ubyte geolocation_flags(time, scanline, ground_pixel) ;
      		geolocation_flags:_FillValue = 255UB ;
      		geolocation_flags:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		geolocation_flags:flag_masks = 0UB, 1UB, 2UB, 4UB, 8UB, 16UB, 32UB, 128UB ;
      		geolocation_flags:flag_meanings = "no_error solar_eclipse sun_glint_possible descending night geo_boundary_crossing spacecraft_manoeuvre geolocation_error" ;
      		geolocation_flags:flag_values = 0UB, 1UB, 2UB, 4UB, 8UB, 16UB, 32UB, 128UB ;
      		geolocation_flags:long_name = "geolocation flags" ;
      		geolocation_flags:max_val = 254UB ;
      		geolocation_flags:min_val = 0UB ;
      		geolocation_flags:units = "1" ;
      } // group GEOLOCATIONS

    group: DETAILED_RESULTS {
      variables:
      	uint processing_quality_flags(time, scanline, ground_pixel) ;
      		processing_quality_flags:long_name = "Processing quality flags" ;
      		processing_quality_flags:comment = "Flags indicating conditions that affect quality of the retrieval." ;
      		processing_quality_flags:flag_meanings = "success radiance_missing irradiance_missing input_spectrum_missing reflectance_range_error ler_range_error snr_range_error sza_range_error vza_range_error lut_range_error ozone_range_error wavelength_offset_error initialization_error memory_error assertion_error io_error numerical_error lut_error ISRF_error convergence_error cloud_filter_convergence_error max_iteration_convergence_error aot_lower_boundary_convergence_error other_boundary_convergence_error geolocation_error ch4_noscat_zero_error h2o_noscat_zero_error max_optical_thickness_error aerosol_boundary_error boundary_hit_error chi2_error svd_error dfs_error radiative_transfer_error optimal_estimation_error profile_error cloud_error model_error number_of_input_data_points_too_low_error cloud_pressure_spread_too_low_error cloud_too_low_level_error generic_range_error generic_exception input_spectrum_alignment_error abort_error wrong_input_type_error wavelength_calibration_error coregistration_error slant_column_density_error airmass_factor_error vertical_column_density_error signal_to_noise_ratio_error configuration_error key_error saturation_error max_num_outlier_exceeded_error solar_eclipse_filter cloud_filter altitude_consistency_filter altitude_roughness_filter sun_glint_filter mixed_surface_type_filter snow_ice_filter aai_filter cloud_fraction_fresco_filter aai_scene_albedo_filter small_pixel_radiance_std_filter cloud_fraction_viirs_filter cirrus_reflectance_viirs_filter cf_viirs_swir_ifov_filter cf_viirs_swir_ofova_filter cf_viirs_swir_ofovb_filter cf_viirs_swir_ofovc_filter cf_viirs_nir_ifov_filter cf_viirs_nir_ofova_filter cf_viirs_nir_ofovb_filter cf_viirs_nir_ofovc_filter refl_cirrus_viirs_swir_filter refl_cirrus_viirs_nir_filter diff_refl_cirrus_viirs_filter ch4_noscat_ratio_filter ch4_noscat_ratio_std_filter h2o_noscat_ratio_filter h2o_noscat_ratio_std_filter diff_psurf_fresco_ecmwf_filter psurf_fresco_stdv_filter ocean_filter time_range_filter pixel_or_scanline_index_filter geographic_region_filter internal_cloud_mask_filter input_spectrum_warning wavelength_calibration_warning extrapolation_warning sun_glint_warning south_atlantic_anomaly_warning sun_glint_correction snow_ice_warning cloud_warning AAI_warning pixel_level_input_data_missing data_range_warning low_cloud_fraction_warning altitude_consistency_warning signal_to_noise_ratio_warning deconvolution_warning so2_volcanic_origin_likely_warning so2_volcanic_origin_certain_warning interpolation_warning saturation_warning high_sza_warning cloud_retrieval_warning cloud_inhomogeneity_warning thermal_instability_warning" ;
      		processing_quality_flags:flag_masks = 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 256U, 512U, 1024U, 2048U, 4096U, 8192U, 16384U, 32768U, 65536U, 131072U, 262144U, 524288U, 1048576U, 2097152U, 4194304U, 8388608U, 16777216U, 33554432U, 67108864U, 134217728U, 268435456U, 536870912U, 1073741824U ;
      		processing_quality_flags:flag_values = 0U, 1U, 2U, 3U, 4U, 5U, 6U, 7U, 8U, 9U, 10U, 11U, 12U, 13U, 14U, 15U, 16U, 17U, 18U, 19U, 20U, 21U, 22U, 23U, 24U, 25U, 26U, 27U, 28U, 29U, 30U, 31U, 32U, 33U, 34U, 35U, 36U, 37U, 38U, 39U, 40U, 41U, 42U, 43U, 44U, 45U, 46U, 47U, 48U, 49U, 50U, 51U, 52U, 53U, 54U, 55U, 64U, 65U, 66U, 67U, 68U, 69U, 70U, 71U, 72U, 73U, 74U, 75U, 76U, 77U, 78U, 79U, 80U, 81U, 82U, 83U, 84U, 85U, 86U, 87U, 88U, 89U, 90U, 91U, 92U, 93U, 94U, 95U, 96U, 97U, 98U, 256U, 512U, 1024U, 2048U, 4096U, 8192U, 16384U, 32768U, 65536U, 131072U, 262144U, 524288U, 1048576U, 2097152U, 4194304U, 8388608U, 16777216U, 33554432U, 67108864U, 134217728U, 268435456U, 536870912U, 1073741824U ;
      		processing_quality_flags:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		processing_quality_flags:_FillValue = 4294967295U ;
      	ushort number_of_spectral_points_in_retrieval(time, scanline, ground_pixel) ;
      		number_of_spectral_points_in_retrieval:long_name = "Number of spectral points used in the retrieval" ;
      		number_of_spectral_points_in_retrieval:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		number_of_spectral_points_in_retrieval:_FillValue = 65535US ;
      	ushort number_of_spectral_points_in_retrieval_NIR(time, scanline, ground_pixel) ;
      		number_of_spectral_points_in_retrieval_NIR:long_name = "number of spectral points used in the retrieval." ;
      		number_of_spectral_points_in_retrieval_NIR:comment = "Flags indicating conditions that affect quality of the retrieval." ;
      		number_of_spectral_points_in_retrieval_NIR:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		number_of_spectral_points_in_retrieval_NIR:_FillValue = 65535US ;
      	float column_averaging_kernel(time, scanline, ground_pixel, layer) ;
      		column_averaging_kernel:units = "1" ;
      		column_averaging_kernel:long_name = "Column averaging kernel for the methane retrieval" ;
      		column_averaging_kernel:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		column_averaging_kernel:_FillValue = 9.96921e+36f ;
      	float carbonmonoxide_total_column(time, scanline, ground_pixel) ;
      		carbonmonoxide_total_column:units = "mol m-2" ;
      		carbonmonoxide_total_column:standard_name = "atmosphere_mole_content_of_carbon_monoxide" ;
      		carbonmonoxide_total_column:long_name = "CO total vertical column" ;
      		carbonmonoxide_total_column:comment = "This is a by-product of the methane retrieval, this is not the official carbon monoxide product." ;
      		carbonmonoxide_total_column:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		carbonmonoxide_total_column:multiplication_factor_to_convert_to_molecules_percm2 = 6.022141e+19f ;
      		carbonmonoxide_total_column:_FillValue = 9.96921e+36f ;
      	float carbonmonoxide_total_column_precision(time, scanline, ground_pixel) ;
      		carbonmonoxide_total_column_precision:units = "mol m-2" ;
      		carbonmonoxide_total_column_precision:standard_name = "atmosphere_mole_content_of_carbon_monoxide standard_error" ;
      		carbonmonoxide_total_column_precision:long_name = "CO total vertical column precision" ;
      		carbonmonoxide_total_column_precision:comment = "This is a by-product of the methane retrieval, this is not the official carbon monoxide product." ;
      		carbonmonoxide_total_column_precision:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		carbonmonoxide_total_column_precision:multiplication_factor_to_convert_to_molecules_percm2 = 6.022141e+19f ;
      		carbonmonoxide_total_column_precision:_FillValue = 9.96921e+36f ;
      	float water_total_column(time, scanline, ground_pixel) ;
      		water_total_column:units = "mol m-2" ;
      		water_total_column:standard_name = "atmosphere_mole_content_of_water_vapor" ;
      		water_total_column:long_name = "H2O total vertical column" ;
      		water_total_column:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		water_total_column:multiplication_factor_to_convert_to_molecules_percm2 = 6.022141e+19f ;
      		water_total_column:_FillValue = 9.96921e+36f ;
      	float water_total_column_precision(time, scanline, ground_pixel) ;
      		water_total_column_precision:units = "mol m-2" ;
      		water_total_column_precision:standard_name = "atmosphere_mole_content_of_water_vapor standard_error" ;
      		water_total_column_precision:long_name = "H2O total vertical column precision" ;
      		water_total_column_precision:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		water_total_column_precision:multiplication_factor_to_convert_to_molecules_percm2 = 6.022141e+19f ;
      		water_total_column_precision:_FillValue = 9.96921e+36f ;
      	float aerosol_size(time, scanline, ground_pixel) ;
      		aerosol_size:units = "1" ;
      		aerosol_size:long_name = "aerosol size parameter of the power law size distribution" ;
      		aerosol_size:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		aerosol_size:_FillValue = 9.96921e+36f ;
      	float aerosol_size_precision(time, scanline, ground_pixel) ;
      		aerosol_size_precision:units = "1" ;
      		aerosol_size_precision:long_name = "precision of the aerosol size parameter of the power law size distribution" ;
      		aerosol_size_precision:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		aerosol_size_precision:_FillValue = 9.96921e+36f ;
      	float aerosol_number_column(time, scanline, ground_pixel) ;
      		aerosol_number_column:units = "m-2" ;
      		aerosol_number_column:standard_name = "atmosphere_number_content_of_aerosol_particles" ;
      		aerosol_number_column:long_name = "aerosol total vertical number column" ;
      		aerosol_number_column:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		aerosol_number_column:_FillValue = 9.96921e+36f ;
      	float aerosol_number_column_precision(time, scanline, ground_pixel) ;
      		aerosol_number_column_precision:units = "m-2" ;
      		aerosol_number_column_precision:standard_name = "atmosphere_number_content_of_aerosol_particles standard_error" ;
      		aerosol_number_column_precision:long_name = "precision of aerosol total vertical column" ;
      		aerosol_number_column_precision:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		aerosol_number_column_precision:_FillValue = 9.96921e+36f ;
      	float aerosol_mid_altitude(time, scanline, ground_pixel) ;
      		aerosol_mid_altitude:units = "m" ;
      		aerosol_mid_altitude:long_name = "central altitude of aerosol altitude distribution. This is the geometric height above the geoid." ;
      		aerosol_mid_altitude:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		aerosol_mid_altitude:_FillValue = 9.96921e+36f ;
      	float aerosol_mid_altitude_precision(time, scanline, ground_pixel) ;
      		aerosol_mid_altitude_precision:units = "m" ;
      		aerosol_mid_altitude_precision:long_name = "precision of central altitude of aerosol altitude distribution." ;
      		aerosol_mid_altitude_precision:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		aerosol_mid_altitude_precision:_FillValue = 9.96921e+36f ;
      	float surface_albedo_SWIR(time, scanline, ground_pixel) ;
      		surface_albedo_SWIR:units = "1" ;
      		surface_albedo_SWIR:standard_name = "surface_albedo" ;
      		surface_albedo_SWIR:long_name = "surface albedo in the SWIR channel" ;
      		surface_albedo_SWIR:radiation_wavelength = 2345.f ;
      		surface_albedo_SWIR:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		surface_albedo_SWIR:_FillValue = 9.96921e+36f ;
      	float surface_albedo_SWIR_precision(time, scanline, ground_pixel) ;
      		surface_albedo_SWIR_precision:units = "1" ;
      		surface_albedo_SWIR_precision:standard_name = "surface_albedo standard_error" ;
      		surface_albedo_SWIR_precision:long_name = "precision of the surface albedo in the SWIR channel" ;
      		surface_albedo_SWIR_precision:radiation_wavelength = 2345.f ;
      		surface_albedo_SWIR_precision:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		surface_albedo_SWIR_precision:_FillValue = 9.96921e+36f ;
      	float surface_albedo_NIR(time, scanline, ground_pixel) ;
      		surface_albedo_NIR:units = "1" ;
      		surface_albedo_NIR:standard_name = "surface_albedo" ;
      		surface_albedo_NIR:long_name = "surface albedo in the NIR channel" ;
      		surface_albedo_NIR:radiation_wavelength = 758.f ;
      		surface_albedo_NIR:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		surface_albedo_NIR:_FillValue = 9.96921e+36f ;
      	float surface_albedo_NIR_precision(time, scanline, ground_pixel) ;
      		surface_albedo_NIR_precision:units = "1" ;
      		surface_albedo_NIR_precision:standard_name = "surface_albedo standard_error" ;
      		surface_albedo_NIR_precision:long_name = "precision of the surface albedo in the NIR channel" ;
      		surface_albedo_NIR_precision:radiation_wavelength = 758.f ;
      		surface_albedo_NIR_precision:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		surface_albedo_NIR_precision:_FillValue = 9.96921e+36f ;
      	float aerosol_optical_thickness_SWIR(time, scanline, ground_pixel) ;
      		aerosol_optical_thickness_SWIR:units = "1" ;
      		aerosol_optical_thickness_SWIR:long_name = "aerosol optical thickness in SWIR channel" ;
      		aerosol_optical_thickness_SWIR:radiation_wavelength = 2345.f ;
      		aerosol_optical_thickness_SWIR:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		aerosol_optical_thickness_SWIR:_FillValue = 9.96921e+36f ;
      	float aerosol_optical_thickness_NIR(time, scanline, ground_pixel) ;
      		aerosol_optical_thickness_NIR:units = "1" ;
      		aerosol_optical_thickness_NIR:long_name = "aerosol optical thickness in NIR band" ;
      		aerosol_optical_thickness_NIR:radiation_wavelength = 758.f ;
      		aerosol_optical_thickness_NIR:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		aerosol_optical_thickness_NIR:_FillValue = 9.96921e+36f ;
      	float wavelength_calibration_offset_SWIR(time, scanline, ground_pixel) ;
      		wavelength_calibration_offset_SWIR:units = "nm" ;
      		wavelength_calibration_offset_SWIR:long_name = "Spectral shift in the SWIR band, add value to L1B to obtain best fit result" ;
      		wavelength_calibration_offset_SWIR:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		wavelength_calibration_offset_SWIR:_FillValue = 9.96921e+36f ;
      	float wavelength_calibration_offset_NIR(time, scanline, ground_pixel) ;
      		wavelength_calibration_offset_NIR:units = "nm" ;
      		wavelength_calibration_offset_NIR:long_name = "Spectral shift in the NIR band, add value to L1B to obtain best fit result" ;
      		wavelength_calibration_offset_NIR:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		wavelength_calibration_offset_NIR:_FillValue = 9.96921e+36f ;
      	float maximum_reflectance_NIR(time, scanline, ground_pixel) ;
      		maximum_reflectance_NIR:units = "1" ;
      		maximum_reflectance_NIR:long_name = "Maximum reflectance in the NIR channel" ;
      		maximum_reflectance_NIR:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		maximum_reflectance_NIR:_FillValue = 9.96921e+36f ;
      	float maximum_reflectance_SWIR(time, scanline, ground_pixel) ;
      		maximum_reflectance_SWIR:units = "1" ;
      		maximum_reflectance_SWIR:long_name = "Maximum reflectance in the SWIR channel" ;
      		maximum_reflectance_SWIR:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		maximum_reflectance_SWIR:_FillValue = 9.96921e+36f ;
      	float chi_square(time, scanline, ground_pixel) ;
      		chi_square:units = "1" ;
      		chi_square:long_name = "chi squared of fit in both SWIR and NIR band" ;
      		chi_square:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		chi_square:_FillValue = 9.96921e+36f ;
      	float chi_square_SWIR(time, scanline, ground_pixel) ;
      		chi_square_SWIR:units = "1" ;
      		chi_square_SWIR:long_name = "chi squared of fit in SWIR band" ;
      		chi_square_SWIR:radiation_wavelength = 2345.f ;
      		chi_square_SWIR:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		chi_square_SWIR:_FillValue = 9.96921e+36f ;
      	float chi_square_NIR(time, scanline, ground_pixel) ;
      		chi_square_NIR:units = "1" ;
      		chi_square_NIR:long_name = "chi squared of fit in NIR band" ;
      		chi_square_NIR:radiation_wavelength = 758.f ;
      		chi_square_NIR:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		chi_square_NIR:_FillValue = 9.96921e+36f ;
      	float degrees_of_freedom(time, scanline, ground_pixel) ;
      		degrees_of_freedom:units = "1" ;
      		degrees_of_freedom:long_name = "degrees of freedom for signal" ;
      		degrees_of_freedom:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		degrees_of_freedom:_FillValue = 9.96921e+36f ;
      	float degrees_of_freedom_methane(time, scanline, ground_pixel) ;
      		degrees_of_freedom_methane:units = "1" ;
      		degrees_of_freedom_methane:long_name = "degrees of freedom for \\Methane profile" ;
      		degrees_of_freedom_methane:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		degrees_of_freedom_methane:_FillValue = 9.96921e+36f ;
      	float degrees_of_freedom_aerosol(time, scanline, ground_pixel) ;
      		degrees_of_freedom_aerosol:units = "1" ;
      		degrees_of_freedom_aerosol:long_name = "degrees of freedom for aerosol parameters" ;
      		degrees_of_freedom_aerosol:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		degrees_of_freedom_aerosol:_FillValue = 9.96921e+36f ;
      	int number_of_iterations(time, scanline, ground_pixel) ;
      		number_of_iterations:long_name = "number of iterations" ;
      		number_of_iterations:units = "1" ;
      		number_of_iterations:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		number_of_iterations:_FillValue = -2147483647 ;
      	float fluorescence(time, scanline, ground_pixel) ;
      		fluorescence:units = "mol s-1 m-2 nm-1 sr-1" ;
      		fluorescence:long_name = "fluorescence emission" ;
      		fluorescence:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		fluorescence:multiplication_factor_to_convert_to_photons_persecond_pernm_percm2_persr = 6.022141e+19f ;
      		fluorescence:_FillValue = 9.96921e+36f ;
      } // group DETAILED_RESULTS

    group: INPUT_DATA {
      variables:
      	float surface_altitude(time, scanline, ground_pixel) ;
      		surface_altitude:long_name = "Surface altitude" ;
      		surface_altitude:standard_name = "surface_altitude" ;
      		surface_altitude:units = "m" ;
      		surface_altitude:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		surface_altitude:source = "http://topotools.cr.usgs.gov/gmted_viewer/" ;
      		surface_altitude:comment = "The mean of the sub-pixels of the surface altitudewithin the approximate field of view, based on the GMTED2010 surface elevation database" ;
      		surface_altitude:_FillValue = 9.96921e+36f ;
      	float surface_altitude_precision(time, scanline, ground_pixel) ;
      		surface_altitude_precision:long_name = "surface altitude precision" ;
      		surface_altitude_precision:standard_name = "surface_altitude standard_error" ;
      		surface_altitude_precision:units = "m" ;
      		surface_altitude_precision:standard_error_multiplier = 1.f ;
      		surface_altitude_precision:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		surface_altitude_precision:source = "http://topotools.cr.usgs.gov/gmted_viewer/" ;
      		surface_altitude_precision:comment = "The standard deviation of sub-pixels used in calculating the mean surface altitude, based on the GMTED2010 surface elevation database" ;
      		surface_altitude_precision:_FillValue = 9.96921e+36f ;
      	ubyte surface_classification(time, scanline, ground_pixel) ;
      		surface_classification:long_name = "Land-water mask and surface classification based on a static database" ;
      		surface_classification:comment = "Flag indicating land/water and further surface classifications for the ground pixel" ;
      		surface_classification:source = "USGS (https://lta.cr.usgs.gov/GLCC) and NASA SDP toolkit (http://newsroom.gsfc.nasa.gov/sdptoolkit/toolkit.html)" ;
      		surface_classification:flag_meanings = "land water some_water coast value_covers_majority_of_pixel water+shallow_ocean water+shallow_inland_water water+ocean_coastline-lake_shoreline water+intermittent_water water+deep_inland_water water+continental_shelf_ocean water+deep_ocean land+urban_and_built-up_land land+dryland_cropland_and_pasture land+irrigated_cropland_and_pasture land+mixed_dryland-irrigated_cropland_and_pasture land+cropland-grassland_mosaic land+cropland-woodland_mosaic land+grassland land+shrubland land+mixed_shrubland-grassland land+savanna land+deciduous_broadleaf_forest land+deciduous_needleleaf_forest land+evergreen_broadleaf_forest land+evergreen_needleleaf_forest land+mixed_forest land+herbaceous_wetland land+wooded_wetland land+barren_or_sparsely_vegetated land+herbaceous_tundra land+wooded_tundra land+mixed_tundra land+bare_ground_tundra land+snow_or_ice" ;
      		surface_classification:flag_values = 0UB, 1UB, 2UB, 3UB, 4UB, 9UB, 17UB, 25UB, 33UB, 41UB, 49UB, 57UB, 8UB, 16UB, 24UB, 32UB, 40UB, 48UB, 56UB, 64UB, 72UB, 80UB, 88UB, 96UB, 104UB, 112UB, 120UB, 128UB, 136UB, 144UB, 152UB, 160UB, 168UB, 176UB, 184UB ;
      		surface_classification:flag_masks = 3UB, 3UB, 3UB, 3UB, 4UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB ;
      		surface_classification:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		surface_classification:_FillValue = 255UB ;
      	int instrument_configuration_identifier(time, scanline) ;
      		instrument_configuration_identifier:long_name = "IcID" ;
      		instrument_configuration_identifier:comment = "The Instrument Configuration ID defines the type of measurement and its purpose. The number of instrument configuration IDs will increase over the mission as new types of measurements are created and used" ;
      		instrument_configuration_identifier:_FillValue = -2147483647 ;
      	short instrument_configuration_version(time, scanline) ;
      		instrument_configuration_version:long_name = "IcVersion" ;
      		instrument_configuration_version:comment = "Version of the instrument_configuration_identifier" ;
      		instrument_configuration_version:_FillValue = -32767s ;
      	float scaled_small_pixel_variance(time, scanline, ground_pixel) ;
      		scaled_small_pixel_variance:long_name = "scaled small pixel variance" ;
      		scaled_small_pixel_variance:units = "1" ;
      		scaled_small_pixel_variance:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		scaled_small_pixel_variance:comment = "The scaled variance of the reflectances of the small pixels" ;
      		scaled_small_pixel_variance:radiation_wavelength = 2315.f ;
      		scaled_small_pixel_variance:_FillValue = 9.96921e+36f ;
      	float eastward_wind(time, scanline, ground_pixel) ;
      		eastward_wind:standard_name = "eastward_wind" ;
      		eastward_wind:long_name = "Eastward wind from ECMWF at 10 meter height level" ;
      		eastward_wind:units = "m s-1" ;
      		eastward_wind:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		eastward_wind:ancillary_variables = "northward_wind" ;
      		eastward_wind:_FillValue = 9.96921e+36f ;
      	float northward_wind(time, scanline, ground_pixel) ;
      		northward_wind:standard_name = "northward_wind" ;
      		northward_wind:long_name = "Northward wind from ECMWF at 10 meter height level" ;
      		northward_wind:units = "m s-1" ;
      		northward_wind:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		northward_wind:ancillary_variables = "eastward_wind" ;
      		northward_wind:_FillValue = 9.96921e+36f ;
      	float methane_profile_apriori(time, scanline, ground_pixel, layer) ;
      		methane_profile_apriori:units = "mol m-2" ;
      		methane_profile_apriori:standard_name = "mole_content_of_methane_in_atmosphere_layer" ;
      		methane_profile_apriori:long_name = "mole content of methane in atmosphere layer" ;
      		methane_profile_apriori:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		methane_profile_apriori:multiplication_factor_to_convert_to_molecules_percm2 = 6.022141e+19f ;
      		methane_profile_apriori:_FillValue = 9.96921e+36f ;
      	float altitude_levels(time, scanline, ground_pixel, level) ;
      		altitude_levels:units = "m" ;
      		altitude_levels:standard_name = "altitude" ;
      		altitude_levels:long_name = "height above the geoid" ;
      		altitude_levels:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		altitude_levels:_FillValue = 9.96921e+36f ;
      	float dry_air_subcolumns(time, scanline, ground_pixel, layer) ;
      		dry_air_subcolumns:units = "mol m-2" ;
      		dry_air_subcolumns:proposed_standard_name = "mole_content_of_dry_air_in_atmosphere_layer" ;
      		dry_air_subcolumns:long_name = "dry air subcolumns" ;
      		dry_air_subcolumns:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		dry_air_subcolumns:multiplication_factor_to_convert_to_molecules_percm2 = 6.022141e+19f ;
      		dry_air_subcolumns:_FillValue = 9.96921e+36f ;
      	float surface_pressure(time, scanline, ground_pixel) ;
      		surface_pressure:units = "Pa" ;
      		surface_pressure:standard_name = "surface_air_pressure" ;
      		surface_pressure:long_name = "surface air pressure" ;
      		surface_pressure:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		surface_pressure:_FillValue = 9.96921e+36f ;
      	float pressure_interval(time, scanline, ground_pixel) ;
      		pressure_interval:units = "Pa" ;
      		pressure_interval:long_name = "pressure difference between levels in the retrieval" ;
      		pressure_interval:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		pressure_interval:_FillValue = 9.96921e+36f ;
      	float cloud_fraction_VIIRS_SWIR_IFOV(time, scanline, ground_pixel) ;
      		cloud_fraction_VIIRS_SWIR_IFOV:units = "1" ;
      		cloud_fraction_VIIRS_SWIR_IFOV:long_name = "Cloud fraction from VIIRS data in the SWIR channel for the instantaneous field of view" ;
      		cloud_fraction_VIIRS_SWIR_IFOV:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		cloud_fraction_VIIRS_SWIR_IFOV:_FillValue = 9.96921e+36f ;
      	float cloud_fraction_VIIRS_SWIR_OFOVa(time, scanline, ground_pixel) ;
      		cloud_fraction_VIIRS_SWIR_OFOVa:units = "1" ;
      		cloud_fraction_VIIRS_SWIR_OFOVa:long_name = "Cloud fraction from VIIRS data in the SWIR channel for the 10% upscaled field of view" ;
      		cloud_fraction_VIIRS_SWIR_OFOVa:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		cloud_fraction_VIIRS_SWIR_OFOVa:_FillValue = 9.96921e+36f ;
      	float cloud_fraction_VIIRS_SWIR_OFOVb(time, scanline, ground_pixel) ;
      		cloud_fraction_VIIRS_SWIR_OFOVb:units = "1" ;
      		cloud_fraction_VIIRS_SWIR_OFOVb:long_name = "Cloud fraction from VIIRS data in the SWIR channel for the 50% upscaled field of view" ;
      		cloud_fraction_VIIRS_SWIR_OFOVb:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		cloud_fraction_VIIRS_SWIR_OFOVb:_FillValue = 9.96921e+36f ;
      	float cloud_fraction_VIIRS_SWIR_OFOVc(time, scanline, ground_pixel) ;
      		cloud_fraction_VIIRS_SWIR_OFOVc:units = "1" ;
      		cloud_fraction_VIIRS_SWIR_OFOVc:long_name = "Cloud fraction from VIIRS data in the SWIR channel for the 100% upscaled field of view" ;
      		cloud_fraction_VIIRS_SWIR_OFOVc:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		cloud_fraction_VIIRS_SWIR_OFOVc:_FillValue = 9.96921e+36f ;
      	float cloud_fraction_VIIRS_NIR_IFOV(time, scanline, ground_pixel) ;
      		cloud_fraction_VIIRS_NIR_IFOV:units = "1" ;
      		cloud_fraction_VIIRS_NIR_IFOV:long_name = "Cloud fraction from VIIRS data in the NIR channel for the instantaneous field of view (band 6)." ;
      		cloud_fraction_VIIRS_NIR_IFOV:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		cloud_fraction_VIIRS_NIR_IFOV:_FillValue = 9.96921e+36f ;
      	float cloud_fraction_VIIRS_NIR_OFOVa(time, scanline, ground_pixel) ;
      		cloud_fraction_VIIRS_NIR_OFOVa:units = "1" ;
      		cloud_fraction_VIIRS_NIR_OFOVa:long_name = "Cloud fraction from VIIRS data in the SWIR channel for the 10% upscaled field of view" ;
      		cloud_fraction_VIIRS_NIR_OFOVa:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		cloud_fraction_VIIRS_NIR_OFOVa:_FillValue = 9.96921e+36f ;
      	float cloud_fraction_VIIRS_NIR_OFOVb(time, scanline, ground_pixel) ;
      		cloud_fraction_VIIRS_NIR_OFOVb:units = "1" ;
      		cloud_fraction_VIIRS_NIR_OFOVb:long_name = "Cloud fraction from VIIRS data in the SWIR channel for the 50% upscaled field of view" ;
      		cloud_fraction_VIIRS_NIR_OFOVb:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		cloud_fraction_VIIRS_NIR_OFOVb:_FillValue = 9.96921e+36f ;
      	float cloud_fraction_VIIRS_NIR_OFOVc(time, scanline, ground_pixel) ;
      		cloud_fraction_VIIRS_NIR_OFOVc:units = "1" ;
      		cloud_fraction_VIIRS_NIR_OFOVc:long_name = "Cloud fraction from VIIRS data in the SWIR channel for the 100% upscaled field of view" ;
      		cloud_fraction_VIIRS_NIR_OFOVc:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		cloud_fraction_VIIRS_NIR_OFOVc:_FillValue = 9.96921e+36f ;
      	float reflectance_cirrus_VIIRS_SWIR(time, scanline, ground_pixel) ;
      		reflectance_cirrus_VIIRS_SWIR:units = "1" ;
      		reflectance_cirrus_VIIRS_SWIR:long_name = "Cirrus reflectance from VIIRS for the SWIR ground pixel" ;
      		reflectance_cirrus_VIIRS_SWIR:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		reflectance_cirrus_VIIRS_SWIR:_FillValue = 9.96921e+36f ;
      	float reflectance_cirrus_VIIRS_NIR(time, scanline, ground_pixel) ;
      		reflectance_cirrus_VIIRS_NIR:units = "1" ;
      		reflectance_cirrus_VIIRS_NIR:long_name = "Cirrus reflectance from VIIRS for the NIR ground pixel" ;
      		reflectance_cirrus_VIIRS_NIR:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		reflectance_cirrus_VIIRS_NIR:_FillValue = 9.96921e+36f ;
      	ubyte internal_cloud_mask(time, scanline, ground_pixel) ;
      		internal_cloud_mask:units = "1" ;
      		internal_cloud_mask:long_name = "Cloud mask based on CO input data" ;
      		internal_cloud_mask:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		internal_cloud_mask:flag_values = 1UB, 2UB, 4UB, 8UB ;
      		internal_cloud_mask:flag_masks = 1UB, 2UB, 4UB, 8UB ;
      		internal_cloud_mask:flag_meanings = "cloudy_post_1pmlle cloudy_pre_2pct cloudy_pre_10pct prefiltered" ;
      		internal_cloud_mask:comment = "Number of orbits in random forest: 300, 300, 250." ;
      		internal_cloud_mask:_FillValue = 255UB ;
      	float apparent_scene_pressure(time, scanline, ground_pixel) ;
      		apparent_scene_pressure:units = "Pa" ;
      		apparent_scene_pressure:long_name = "Apparent scene pressure from oxygen A-band depth" ;
      		apparent_scene_pressure:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		apparent_scene_pressure:_FillValue = 9.96921e+36f ;
      	float apparent_scene_pressure_standard_deviation(time, scanline, ground_pixel) ;
      		apparent_scene_pressure_standard_deviation:units = "Pa" ;
      		apparent_scene_pressure_standard_deviation:long_name = "Standard deviation of the apparent scene pressure from oxygen A-band depth over 9 ground pixels" ;
      		apparent_scene_pressure_standard_deviation:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		apparent_scene_pressure_standard_deviation:_FillValue = 9.96921e+36f ;
      	float methane_weak_twoband_total_column(time, scanline, ground_pixel) ;
      		methane_weak_twoband_total_column:units = "mol m-2" ;
      		methane_weak_twoband_total_column:standard_name = "atmosphere_mole_content_of_methane" ;
      		methane_weak_twoband_total_column:long_name = "Vertically integrated CH4 column from weak band" ;
      		methane_weak_twoband_total_column:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		methane_weak_twoband_total_column:multiplication_factor_to_convert_to_molecules_percm2 = 6.022141e+19f ;
      		methane_weak_twoband_total_column:_FillValue = 9.96921e+36f ;
      	float methane_strong_twoband_total_column(time, scanline, ground_pixel) ;
      		methane_strong_twoband_total_column:units = "mol m-2" ;
      		methane_strong_twoband_total_column:standard_name = "atmosphere_mole_content_of_methane" ;
      		methane_strong_twoband_total_column:long_name = "Vertically integrated CH4 column from strong band" ;
      		methane_strong_twoband_total_column:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		methane_strong_twoband_total_column:multiplication_factor_to_convert_to_molecules_percm2 = 6.022141e+19f ;
      		methane_strong_twoband_total_column:_FillValue = 9.96921e+36f ;
      	float methane_ratio_weak_strong_standard_deviation(time, scanline, ground_pixel) ;
      		methane_ratio_weak_strong_standard_deviation:units = "1" ;
      		methane_ratio_weak_strong_standard_deviation:long_name = "Standard deviation of ratio of the methane column from weak and strong band over 9 ground pixels" ;
      		methane_ratio_weak_strong_standard_deviation:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		methane_ratio_weak_strong_standard_deviation:_FillValue = 9.96921e+36f ;
      	float water_weak_twoband_total_column(time, scanline, ground_pixel) ;
      		water_weak_twoband_total_column:units = "mol m-2" ;
      		water_weak_twoband_total_column:standard_name = "atmosphere_mole_content_of_water_vapor" ;
      		water_weak_twoband_total_column:long_name = "Vertically integrated H2O column from weak band" ;
      		water_weak_twoband_total_column:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		water_weak_twoband_total_column:multiplication_factor_to_convert_to_molecules_percm2 = 6.022141e+19f ;
      		water_weak_twoband_total_column:_FillValue = 9.96921e+36f ;
      	float water_strong_twoband_total_column(time, scanline, ground_pixel) ;
      		water_strong_twoband_total_column:units = "mol m-2" ;
      		water_strong_twoband_total_column:standard_name = "atmosphere_mole_content_of_water_vapor" ;
      		water_strong_twoband_total_column:long_name = "Vertically integrated H2O column from strong band" ;
      		water_strong_twoband_total_column:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		water_strong_twoband_total_column:multiplication_factor_to_convert_to_molecules_percm2 = 6.022141e+19f ;
      		water_strong_twoband_total_column:_FillValue = 9.96921e+36f ;
      	float water_ratio_weak_strong_standard_deviation(time, scanline, ground_pixel) ;
      		water_ratio_weak_strong_standard_deviation:units = "1" ;
      		water_ratio_weak_strong_standard_deviation:long_name = "Standard deviation of ratio of the water vapor column from weak and strong band over 9 ground pixels" ;
      		water_ratio_weak_strong_standard_deviation:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		water_ratio_weak_strong_standard_deviation:_FillValue = 9.96921e+36f ;
      	float fluorescence_apriori(time, scanline, ground_pixel) ;
      		fluorescence_apriori:units = "mol s-1 m-2 nm-1 sr-1" ;
      		fluorescence_apriori:long_name = "a priori fluorescence emission" ;
      		fluorescence_apriori:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		fluorescence_apriori:multiplication_factor_to_convert_to_photons_persecond_pernm_percm2_persr = 6.022141e+19f ;
      		fluorescence_apriori:_FillValue = 9.96921e+36f ;
      } // group INPUT_DATA
    } // group SUPPORT_DATA
  } // group PRODUCT

group: METADATA {

  group: QA_STATISTICS {
    dimensions:
    	vertices = 2 ;
    	XCH4_histogram_axis = 100 ;
    	XCH4_pdf_axis = 400 ;
    variables:
    	float methane_mixing_ratio_histogram_axis(XCH4_histogram_axis) ;
    		methane_mixing_ratio_histogram_axis:units = "1" ;
    		methane_mixing_ratio_histogram_axis:comment = "Histogram axis of methane mixing ratio" ;
    		methane_mixing_ratio_histogram_axis:long_name = "Histogram of the methane mixing ratio" ;
    		methane_mixing_ratio_histogram_axis:bounds = "XCH4_histogram_bounds" ;
    		methane_mixing_ratio_histogram_axis:_FillValue = 9.96921e+36f ;
    	float methane_mixing_ratio_pdf_axis(XCH4_pdf_axis) ;
    		methane_mixing_ratio_pdf_axis:units = "1" ;
    		methane_mixing_ratio_pdf_axis:comment = "Probability density function of methane dry air mixing ratio" ;
    		methane_mixing_ratio_pdf_axis:long_name = "Probability density function of methane dry air mixing ratio" ;
    		methane_mixing_ratio_pdf_axis:bounds = "XCH4_pdf_bounds" ;
    		methane_mixing_ratio_pdf_axis:_FillValue = 9.96921e+36f ;
    	float methane_mixing_ratio_histogram_bounds(XCH4_histogram_axis, vertices) ;
    		methane_mixing_ratio_histogram_bounds:_FillValue = 9.96921e+36f ;
    	float methane_mixing_ratio_pdf_bounds(XCH4_pdf_axis, vertices) ;
    		methane_mixing_ratio_pdf_bounds:_FillValue = 9.96921e+36f ;
    	int methane_mixing_ratio_histogram(XCH4_histogram_axis) ;
    		methane_mixing_ratio_histogram:comment = "Histogram of the Methane dry air mixing ratio" ;
    		methane_mixing_ratio_histogram:number_of_overflow_values = 17 ;
    		methane_mixing_ratio_histogram:number_of_underflow_values = 0 ;
    		methane_mixing_ratio_histogram:_FillValue = -2147483647 ;
    	float methane_mixing_ratio_pdf(XCH4_pdf_axis) ;
    		methane_mixing_ratio_pdf:comment = "Probability density function of the Methane dry air mixing ratio" ;
    		methane_mixing_ratio_pdf:geolocation_sampling_total = 48752.89f ;
    		methane_mixing_ratio_pdf:_FillValue = 9.96921e+36f ;

    // group attributes:
    		:number_of_groundpixels = 803025 ;
    		:number_of_processed_pixels = 803025 ;
    		:number_of_successfully_processed_pixels = 56583 ;
    		:number_of_rejected_pixels_not_enough_spectrum = 0 ;
    		:number_of_failed_retrievals = 746442 ;
    		:number_of_ground_pixels_with_warnings = 90564 ;
    		:number_of_missing_scanlines = 0 ;
    		:number_of_radiance_missing_occurrences = 0 ;
    		:number_of_irradiance_missing_occurrences = 0 ;
    		:number_of_input_spectrum_missing_occurrences = 0 ;
    		:number_of_reflectance_range_error_occurrences = 0 ;
    		:number_of_ler_range_error_occurrences = 0 ;
    		:number_of_snr_range_error_occurrences = 74 ;
    		:number_of_sza_range_error_occurrences = 104331 ;
    		:number_of_vza_range_error_occurrences = 16134 ;
    		:number_of_lut_range_error_occurrences = 0 ;
    		:number_of_ozone_range_error_occurrences = 0 ;
    		:number_of_wavelength_offset_error_occurrences = 0 ;
    		:number_of_initialization_error_occurrences = 0 ;
    		:number_of_memory_error_occurrences = 0 ;
    		:number_of_assertion_error_occurrences = 0 ;
    		:number_of_io_error_occurrences = 0 ;
    		:number_of_numerical_error_occurrences = 0 ;
    		:number_of_lut_error_occurrences = 0 ;
    		:number_of_ISRF_error_occurrences = 0 ;
    		:number_of_convergence_error_occurrences = 2964 ;
    		:number_of_cloud_filter_convergence_error_occurrences = 0 ;
    		:number_of_max_iteration_convergence_error_occurrences = 2 ;
    		:number_of_aot_lower_boundary_convergence_error_occurrences = 0 ;
    		:number_of_other_boundary_convergence_error_occurrences = 0 ;
    		:number_of_geolocation_error_occurrences = 0 ;
    		:number_of_ch4_noscat_zero_error_occurrences = 0 ;
    		:number_of_h2o_noscat_zero_error_occurrences = 0 ;
    		:number_of_max_optical_thickness_error_occurrences = 419 ;
    		:number_of_aerosol_boundary_error_occurrences = 1 ;
    		:number_of_boundary_hit_error_occurrences = 43 ;
    		:number_of_chi2_error_occurrences = 1258 ;
    		:number_of_svd_error_occurrences = 5 ;
    		:number_of_dfs_error_occurrences = 0 ;
    		:number_of_radiative_transfer_error_occurrences = 0 ;
    		:number_of_optimal_estimation_error_occurrences = 0 ;
    		:number_of_profile_error_occurrences = 0 ;
    		:number_of_cloud_error_occurrences = 0 ;
    		:number_of_model_error_occurrences = 0 ;
    		:number_of_number_of_input_data_points_too_low_error_occurrences = 0 ;
    		:number_of_cloud_pressure_spread_too_low_error_occurrences = 0 ;
    		:number_of_cloud_too_low_level_error_occurrences = 0 ;
    		:number_of_generic_range_error_occurrences = 0 ;
    		:number_of_generic_exception_occurrences = 0 ;
    		:number_of_input_spectrum_alignment_error_occurrences = 0 ;
    		:number_of_abort_error_occurrences = 0 ;
    		:number_of_wrong_input_type_error_occurrences = 0 ;
    		:number_of_wavelength_calibration_error_occurrences = 0 ;
    		:number_of_coregistration_error_occurrences = 0 ;
    		:number_of_slant_column_density_error_occurrences = 0 ;
    		:number_of_airmass_factor_error_occurrences = 0 ;
    		:number_of_vertical_column_density_error_occurrences = 0 ;
    		:number_of_signal_to_noise_ratio_error_occurrences = 0 ;
    		:number_of_configuration_error_occurrences = 0 ;
    		:number_of_key_error_occurrences = 0 ;
    		:number_of_saturation_error_occurrences = 0 ;
    		:number_of_max_num_outlier_exceeded_error_occurrences = 0 ;
    		:number_of_solar_eclipse_filter_occurrences = 0 ;
    		:number_of_cloud_filter_occurrences = 0 ;
    		:number_of_altitude_consistency_filter_occurrences = 0 ;
    		:number_of_altitude_roughness_filter_occurrences = 2127 ;
    		:number_of_sun_glint_filter_occurrences = 0 ;
    		:number_of_mixed_surface_type_filter_occurrences = 0 ;
    		:number_of_snow_ice_filter_occurrences = 0 ;
    		:number_of_aai_filter_occurrences = 0 ;
    		:number_of_cloud_fraction_fresco_filter_occurrences = 0 ;
    		:number_of_aai_scene_albedo_filter_occurrences = 0 ;
    		:number_of_small_pixel_radiance_std_filter_occurrences = 0 ;
    		:number_of_cloud_fraction_viirs_filter_occurrences = 0 ;
    		:number_of_cirrus_reflectance_viirs_filter_occurrences = 0 ;
    		:number_of_cf_viirs_swir_ifov_filter_occurrences = 132352 ;
    		:number_of_cf_viirs_swir_ofova_filter_occurrences = 0 ;
    		:number_of_cf_viirs_swir_ofovb_filter_occurrences = 0 ;
    		:number_of_cf_viirs_swir_ofovc_filter_occurrences = 0 ;
    		:number_of_cf_viirs_nir_ifov_filter_occurrences = 0 ;
    		:number_of_cf_viirs_nir_ofova_filter_occurrences = 0 ;
    		:number_of_cf_viirs_nir_ofovb_filter_occurrences = 0 ;
    		:number_of_cf_viirs_nir_ofovc_filter_occurrences = 0 ;
    		:number_of_refl_cirrus_viirs_swir_filter_occurrences = 0 ;
    		:number_of_refl_cirrus_viirs_nir_filter_occurrences = 0 ;
    		:number_of_diff_refl_cirrus_viirs_filter_occurrences = 0 ;
    		:number_of_ch4_noscat_ratio_filter_occurrences = 0 ;
    		:number_of_ch4_noscat_ratio_std_filter_occurrences = 0 ;
    		:number_of_h2o_noscat_ratio_filter_occurrences = 0 ;
    		:number_of_h2o_noscat_ratio_std_filter_occurrences = 0 ;
    		:number_of_diff_psurf_fresco_ecmwf_filter_occurrences = 0 ;
    		:number_of_psurf_fresco_stdv_filter_occurrences = 0 ;
    		:number_of_ocean_filter_occurrences = 486732 ;
    		:number_of_time_range_filter_occurrences = 0 ;
    		:number_of_pixel_or_scanline_index_filter_occurrences = 0 ;
    		:number_of_geographic_region_filter_occurrences = 0 ;
    		:number_of_internal_cloud_mask_filter_occurrences = 0 ;
    		:number_of_input_spectrum_warning_occurrences = 0 ;
    		:number_of_wavelength_calibration_warning_occurrences = 0 ;
    		:number_of_extrapolation_warning_occurrences = 0 ;
    		:number_of_sun_glint_warning_occurrences = 47853 ;
    		:number_of_south_atlantic_anomaly_warning_occurrences = 0 ;
    		:number_of_sun_glint_correction_occurrences = 0 ;
    		:number_of_snow_ice_warning_occurrences = 0 ;
    		:number_of_cloud_warning_occurrences = 17684 ;
    		:number_of_AAI_warning_occurrences = 0 ;
    		:number_of_pixel_level_input_data_missing_occurrences = 0 ;
    		:number_of_data_range_warning_occurrences = 44762 ;
    		:number_of_low_cloud_fraction_warning_occurrences = 0 ;
    		:number_of_altitude_consistency_warning_occurrences = 904 ;
    		:number_of_signal_to_noise_ratio_warning_occurrences = 0 ;
    		:number_of_deconvolution_warning_occurrences = 0 ;
    		:number_of_so2_volcanic_origin_likely_warning_occurrences = 0 ;
    		:number_of_so2_volcanic_origin_certain_warning_occurrences = 0 ;
    		:number_of_interpolation_warning_occurrences = 0 ;
    		:number_of_saturation_warning_occurrences = 0 ;
    		:number_of_high_sza_warning_occurrences = 0 ;
    		:number_of_cloud_retrieval_warning_occurrences = 0 ;
    		:number_of_cloud_inhomogeneity_warning_occurrences = 0 ;
    		:number_of_thermal_instability_warning_occurrences = 0 ;
    		:global_processing_warnings = "None" ;
    		:time_for_algorithm_initialization = 56.574341 ;
    		:time_for_processing = 27688.735877 ;
    		:time_per_pixel = 3.76196148661263 ;
    		:time_standard_deviation_per_pixel = 0.00237292179501523 ;
    } // group QA_STATISTICS

  group: ALGORITHM_SETTINGS {

    // group attributes:
    		:configuration.version.algorithm = "1.6.0" ;
    		:configuration.version.framework = "1.2.0" ;
    		:coregistration.fraction.minimum = "0.0" ;
    		:input.1.band = "7" ;
    		:input.1.irrType = "L1B_IR_SIR" ;
    		:input.1.type = "L1B_RA_BD7" ;
    		:input.2.band = "8" ;
    		:input.2.irrType = "L1B_IR_SIR" ;
    		:input.2.type = "L1B_RA_BD8" ;
    		:input.3.band = "6" ;
    		:input.3.irrType = "L1B_IR_UVN" ;
    		:input.3.type = "L1B_RA_BD6" ;
    		:input.4.band = "7" ;
    		:input.4.type = "L2__CO____" ;
    		:input.5.band = "6" ;
    		:input.5.type = "L2__FRESCO" ;
    		:input.6.band = "6" ;
    		:input.6.required = "false" ;
    		:input.6.type = "L2__NP_BD6" ;
    		:input.7.band = "7" ;
    		:input.7.required = "false" ;
    		:input.7.type = "L2__NP_BD7" ;
    		:input.8.band = "7" ;
    		:input.8.required = "false" ;
    		:input.8.type = "L2__CH4CLD" ;
    		:input.coadd.count = "1" ;
    		:input.count = "8" ;
    		:output.1.band = "7" ;
    		:output.1.config = "cfg/product/product.CH4___.xml" ;
    		:output.1.type = "L2__CH4___" ;
    		:output.compressionLevel = "3" ;
    		:output.count = "1" ;
    		:output.histogram.methane_mixing_ratio.range = "1200, 2000" ;
    		:output.useCompression = "true" ;
    		:output.useFletcher32 = "true" ;
    		:output.useShuffleFilter = "true" ;
    		:processing.algorithm = "CH4___" ;
    		:processing.cirrusReflectanceIndex = "0" ;
    		:processing.correct_surface_pressure_for_altitude = "false" ;
    		:processing.groupDem = "DEM_RADIUS_05000" ;
    		:processing.radianceFractionMinError = "0" ;
    		:processing.radiancePixelsMinError = "0" ;
    		:processing.sgaLimit = "30.0" ;
    		:processing.szaMax = "180.0" ;
    		:processing.szaMin = "0.0" ;
    		:processing.threadStackSize = "50000000" ;
    		:processing.vzaMax = "180.0" ;
    		:processing.vzaMin = "0.0" ;
    		:qa_value.AAI_warning = "100.0" ;
    		:qa_value.altitude_consistency_warning = "100.0" ;
    		:qa_value.cloud_inhomogeneity_warning = "100.0" ;
    		:qa_value.cloud_retrieval_warning = "100.0" ;
    		:qa_value.cloud_warning = "100.0" ;
    		:qa_value.data_range_warning = "40.0" ;
    		:qa_value.deconvolution_warning = "80.0" ;
    		:qa_value.extrapolation_warning = "100.0" ;
    		:qa_value.high_sza_warning = "100.0" ;
    		:qa_value.input_spectrum_warning = "100.0" ;
    		:qa_value.interpolation_warning = "100.0" ;
    		:qa_value.low_cloud_fraction_warning = "90.0" ;
    		:qa_value.pixel_level_input_data_missing = "40.0" ;
    		:qa_value.saturation_warning = "100.0" ;
    		:qa_value.signal_to_noise_ratio_warning = "100.0" ;
    		:qa_value.snow_ice_warning = "100.0" ;
    		:qa_value.so2_volcanic_origin_certain_warning = "100.0" ;
    		:qa_value.so2_volcanic_origin_likely_warning = "100.0" ;
    		:qa_value.south_atlantic_anomaly_warning = "100.0" ;
    		:qa_value.sun_glint_correction = "100.0" ;
    		:qa_value.sun_glint_warning = "100.0" ;
    		:qa_value.thermal_instability_warning = "40.0" ;
    		:qa_value.wavelength_calibration_warning = "100.0" ;
    		:quality_control.missing_input.max_fraction = "0.25" ;
    		:quality_control.missing_scanlines.max_count = "60" ;
    		:quality_control.missing_scanlines.max_fraction = "0.05" ;
    		:quality_control.qa_value.limit = "0.5" ;
    		:quality_control.success.min_fraction = "0.001" ;
    		:joborder.processing.threads = "9" ;
    } // group ALGORITHM_SETTINGS

  group: GRANULE_DESCRIPTION {

    // group attributes:
    		:GranuleStart = "2024-04-07T13:01:21Z" ;
    		:GranuleEnd = "2024-04-07T13:53:37Z" ;
    		:InstrumentName = "TROPOMI" ;
    		:MissionName = "Sentinel-5 precursor" ;
    		:MissionShortName = "S5P" ;
    		:ProcessLevel = "2" ;
    		:ProcessingCenter = "PDGS-OP" ;
    		:ProcessingNode = "s5p-ops2-off-pn19" ;
    		:ProcessorVersion = "2.6.0" ;
    		:ProductFormatVersion = 10600 ;
    		:ProcessingMode = "Offline" ;
    		:LongitudeOfDaysideNadirEquatorCrossing = 0.671685f ;
    		:CollectionIdentifier = "03" ;
    		:ProductShortName = "L2__CH4___" ;
    } // group GRANULE_DESCRIPTION

  group: ISO_METADATA {

    // group attributes:
    		:gmd\:dateStamp = "2015-10-16" ;
    		:gmd\:fileIdentifier = "urn:ogc:def:EOP:ESA:SENTINEL.S5P_TROP_L2__CH4___" ;
    		:gmd\:hierarchyLevelName = "EO Product Collection" ;
    		:gmd\:metadataStandardName = "ISO 19115-2 Geographic Information - Metadata Part 2 Extensions for imagery and gridded data" ;
    		:gmd\:metadataStandardVersion = "ISO 19115-2:2009(E), S5P profile" ;
    		:objectType = "gmi:MI_Metadata" ;

    group: gmd\:language {

      // group attributes:
      		:codeList = "http://www.loc.gov/standards/iso639-2/" ;
      		:codeListValue = "eng" ;
      		:objectType = "gmd:LanguageCode" ;
      } // group gmd\:language

    group: gmd\:characterSet {

      // group attributes:
      		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#MD_CharacterSetCode" ;
      		:codeListValue = "utf8" ;
      		:objectType = "gmd:MD_CharacterSetCode" ;
      } // group gmd\:characterSet

    group: gmd\:hierarchyLevel {

      // group attributes:
      		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#MD_ScopeCode" ;
      		:codeListValue = "series" ;
      		:objectType = "gmd:MD_ScopeCode" ;
      } // group gmd\:hierarchyLevel

    group: gmd\:contact {

      // group attributes:
      		:gmd\:organisationName = "Copernicus Space Component Data Access System,  ESA, Services Coordinated Interface" ;
      		:objectType = "gmd:CI_ResponsibleParty" ;

      group: gmd\:contactInfo {

        // group attributes:
        		:objectType = "gmd:CI_Contact" ;

        group: gmd\:address {

          // group attributes:
          		:gmd\:electronicMailAddress = "EOSupport@copernicus.esa.int" ;
          		:objectType = "gmd:CI_Address" ;
          } // group gmd\:address
        } // group gmd\:contactInfo

      group: gmd\:role {

        // group attributes:
        		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_RoleCode" ;
        		:codeListValue = "pointOfContact" ;
        		:objectType = "gmd:CI_RoleCode" ;
        } // group gmd\:role
      } // group gmd\:contact

    group: gmd\:identificationInfo {

      // group attributes:
      		:gmd\:abstract = "Dry-air mixing ratio of methane for cloud-free observations with a spatial resolution of 5.5x7.0 km2 observed at about 13:30 local solar time from spectra measured by TROPOMI" ;
      		:gmd\:credit = "The Sentinel 5 Precursor TROPOMI Level 2 products are developed with funding from the European Space Agency (ESA), the Netherlands Space Office (NSO), the Belgian Science Policy Office, the German Aerospace Center (DLR) and the Bayerisches Staatsministerium für Wirtschaft und Medien, Energie und Technologie (StMWi)." ;
      		:gmd\:language = "eng" ;
      		:gmd\:topicCategory = "climatologyMeteorologyAtmosphere" ;
      		:objectType = "gmd:MD_DataIdentification" ;

      group: gmd\:citation {

        // group attributes:
        		:gmd\:title = "TROPOMI/S5P Methane 1-Orbit L2 Swath 5.5x7.0km" ;
        		:objectType = "gmd:CI_Citation" ;

        group: gmd\:date {

          // group attributes:
          		:gmd\:date = "2024-04-09" ;
          		:objectType = "gmd:CI_Date" ;

          group: gmd\:dateType {

            // group attributes:
            		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
            		:codeListValue = "creation" ;
            		:objectType = "gmd:CI_DateTypeCode" ;
            } // group gmd\:dateType
          } // group gmd\:date

        group: gmd\:identifier {

          // group attributes:
          		:gmd\:code = "urn:ogc:def:EOP:ESA:SENTINEL.S5P_TROP_L2__CH4___" ;
          		:objectType = "gmd:MD_Identifier" ;
          } // group gmd\:identifier
        } // group gmd\:citation

      group: gmd\:pointOfContact {

        // group attributes:
        		:gmd\:organisationName = "Copernicus Space Component Data Access System,  ESA, Services Coordinated Interface" ;
        		:objectType = "gmd:CI_ResponsibleParty" ;

        group: gmd\:contactInfo {

          // group attributes:
          		:objectType = "gmd:CI_Contact" ;

          group: gmd\:address {

            // group attributes:
            		:gmd\:electronicMailAddress = "EOSupport@copernicus.esa.int" ;
            		:objectType = "gmd:CI_Address" ;
            } // group gmd\:address
          } // group gmd\:contactInfo

        group: gmd\:role {

          // group attributes:
          		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_RoleCode" ;
          		:codeListValue = "distributor" ;
          		:objectType = "gmd:CI_RoleCode" ;
          } // group gmd\:role
        } // group gmd\:pointOfContact

      group: gmd\:descriptiveKeywords\#1 {

        // group attributes:
        		:gmd\:keyword\#1 = "Atmospheric conditions" ;
        		:objectType = "gmd:MD_Keywords" ;

        group: gmd\:type {

          // group attributes:
          		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#MD_KeywordTypeCode" ;
          		:codeListValue = "theme" ;
          		:objectType = "gmd:MD_KeywordTypeCode" ;
          } // group gmd\:type

        group: gmd\:thesaurusName {

          // group attributes:
          		:gmd\:title = "GEMET - INSPIRE themes, version 1.0" ;
          		:objectType = "gmd:CI_Citation" ;

          group: gmd\:date {

            // group attributes:
            		:gmd\:date = "2008-06-01" ;
            		:objectType = "gmd:CI_Date" ;

            group: gmd\:dateType {

              // group attributes:
              		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
              		:codeListValue = "publication" ;
              		:objectType = "gmd:CI_DateTypeCode" ;
              } // group gmd\:dateType
            } // group gmd\:date
          } // group gmd\:thesaurusName
        } // group gmd\:descriptiveKeywords\#1

      group: gmd\:descriptiveKeywords\#2 {

        // group attributes:
        		:gmd\:keyword\#1 = "atmosphere_mole_fraction_of_methane_in_dry_air" ;
        		:objectType = "gmd:MD_Keywords" ;

        group: gmd\:thesaurusName {

          // group attributes:
          		:gmd\:title = "CF Standard Name Table v65" ;
          		:xlink\:href = "http://cfconventions.org/standard-names.html" ;
          		:objectType = "gmd:CI_Citation" ;

          group: gmd\:date {

            // group attributes:
            		:gmd\:date = "2019-04-09" ;
            		:objectType = "gmd:CI_Date" ;

            group: gmd\:dateType {

              // group attributes:
              		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
              		:codeListValue = "publication" ;
              		:objectType = "gmd:CI_DateTypeCode" ;
              } // group gmd\:dateType
            } // group gmd\:date
          } // group gmd\:thesaurusName
        } // group gmd\:descriptiveKeywords\#2

      group: gmd\:resourceConstraints {

        // group attributes:
        		:gmd\:useLimitation = "no conditions apply" ;
        		:objectType = "gmd:MD_LegalConstraints" ;

        group: gmd\:accessConstraints {

          // group attributes:
          		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#MD_RestrictionCode" ;
          		:codeListValue = "copyright" ;
          		:objectType = "gmd:MD_RestrictionCode" ;
          } // group gmd\:accessConstraints
        } // group gmd\:resourceConstraints

      group: gmd\:spatialRepresentationType {

        // group attributes:
        		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#MD_SpatialRepresentationTypeCode" ;
        		:codeListValue = "grid" ;
        		:objectType = "gmd:MD_SpatialRepresentationTypeCode" ;
        } // group gmd\:spatialRepresentationType

      group: gmd\:characterSet {

        // group attributes:
        		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#MD_CharacterSetCode" ;
        		:codeListValue = "utf8" ;
        		:objectType = "gmd:MD_CharacterSetCode" ;
        } // group gmd\:characterSet

      group: gmd\:extent {

        // group attributes:
        		:objectType = "gmd:EX_Extent" ;

        group: gmd\:geographicElement {

          // group attributes:
          		:gmd\:eastBoundLongitude = 179.9852f ;
          		:gmd\:northBoundLatitude = 89.94537f ;
          		:gmd\:southBoundLatitude = -89.94071f ;
          		:gmd\:westBoundLongitude = -179.9215f ;
          		:gmd\:extentTypeCode = "true" ;
          		:objectType = "gmd:EX_GeographicBoundingBox" ;
          } // group gmd\:geographicElement

        group: gmd\:temporalElement {

          // group attributes:
          		:objectType = "gmd:EX_TemporalExtent" ;

          group: gmd\:extent {

            // group attributes:
            		:gml\:beginPosition = "2024-04-07T13:01:21Z" ;
            		:gml\:endPosition = "2024-04-07T13:53:37Z" ;
            		:objectType = "gml:TimePeriod" ;
            } // group gmd\:extent
          } // group gmd\:temporalElement
        } // group gmd\:extent
      } // group gmd\:identificationInfo

    group: gmd\:dataQualityInfo {

      // group attributes:
      		:objectType = "gmd:DQ_DataQuality" ;

      group: gmd\:scope {

        // group attributes:
        		:objectType = "gmd:DQ_Scope" ;

        group: gmd\:level {

          // group attributes:
          		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#MD_ScopeCode" ;
          		:codeListValue = "dataset" ;
          		:objectType = "gmd:MD_ScopeCode" ;
          } // group gmd\:level
        } // group gmd\:scope

      group: gmd\:report {

        // group attributes:
        		:objectType = "gmd:DQ_DomainConsistency" ;

        group: gmd\:result {

          // group attributes:
          		:objectType = "gmd:DQ_ConformanceResult" ;
          		:gmd\:pass = "true" ;
          		:gmd\:explanation = "INSPIRE Data specification for orthoimagery is not yet officially published so conformity has not yet been evaluated" ;

          group: gmd\:specification {

            // group attributes:
            		:objectType = "gmd:CI_Citation" ;
            		:gmd\:title = "INSPIRE Data Specification on Orthoimagery - Guidelines, version 3.0rc3" ;

            group: gmd\:date {

              // group attributes:
              		:gmd\:date = "2013-02-04" ;
              		:objectType = "gmd:CI_Date" ;

              group: gmd\:dateType {

                // group attributes:
                		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                		:codeListValue = "publication" ;
                		:objectType = "gmd:CI_DateTypeCode" ;
                } // group gmd\:dateType
              } // group gmd\:date
            } // group gmd\:specification
          } // group gmd\:result
        } // group gmd\:report

      group: gmd\:lineage {

        // group attributes:
        		:objectType = "gmd:LI_Lineage" ;
        		:gmd\:statement = "L2 CH4___ dataset produced by PDGS-OP from the S5P/TROPOMI L1B product" ;

        group: gmd\:processStep {

          // group attributes:
          		:objectType = "gmi:LE_ProcessStep" ;
          		:gmd\:description = "Processing of L1b to L2 CH4___ data for orbit 33598 using the KNMI/SRON processor version 2.6.0" ;

          group: gmi\:output {

            // group attributes:
            		:gmd\:description = "TROPOMI/S5P Methane 1-Orbit L2 Swath 5.5x7.0km" ;
            		:objectType = "gmi:LE_Source" ;

            group: gmd\:sourceCitation {

              // group attributes:
              		:gmd\:title = "S5P_OFFL_L2__CH4____20240407T123946_20240407T142117_33598_03_020600_20240409T045638" ;
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2024-04-09" ;
                		:objectType = "gmd:CI_DateTime" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:identifier {

                // group attributes:
                		:gmd\:code = "L2__CH4___" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmd\:identifier
              } // group gmd\:sourceCitation

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "L2" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel
            } // group gmi\:output

          group: gmi\:processingInformation {

            // group attributes:
            		:objectType = "gmi:LE_Processing" ;

            group: gmi\:identifier {

              // group attributes:
              		:gmd\:code = "KNMI/SRON L2 CH4___ processor, version 2.6.0" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:identifier

            group: gmi\:softwareReference {

              // group attributes:
              		:gmd\:title = "TROPNLL2DP processor" ;
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2023-09-28T07:04:00Z" ;
                		:objectType = "gmd:CI_DateTime" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date
              } // group gmi\:softwareReference

            group: gmi\:documentation\#1 {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;
              		:gmd\:title = "Algorithm Theoretical Baseline Document for Sentinel-5 Precursor Methane Retrieval; SRON-S5P-LEV2-RP-001; release 1.0" ;
              		:doi = "N/A" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2015-11-30" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "revision" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date
              } // group gmi\:documentation\#1

            group: gmi\:documentation\#2 {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;
              		:gmd\:title = "Sentinel-5 precursor/TROPOMI Level 2 Product User Manual Methane; SRON-S5P-LEV2-MA-001; release 1.0" ;
              		:doi = "N/A" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2015-11-30" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "revision" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date
              } // group gmi\:documentation\#2
            } // group gmi\:processingInformation

          group: gmi\:report {

            // group attributes:
            		:gmi\:description = "Sentinel 5-precursor TROPOMI L1b processed to L2 data using the KNMI/SRON L2 CH4___ processor" ;
            		:gmi\:fileType = "netCDF-4" ;
            		:gmi\:name = "S5P_OFFL_L2__CH4____20240407T123946_20240407T142117_33598_03_020600_20240409T045638.nc" ;
            		:objectType = "gmi:LE_ProcessStepReport" ;
            } // group gmi\:report

          group: gmd\:source\#1 {

            // group attributes:
            		:objectType = "gmi:LE_Source" ;
            		:gmd\:description = "Auxiliary CTM AUX_CTMCH4 model input data" ;

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "N/A" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2024-04-09T12:47:23Z" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:title {

                // group attributes:
                		:gco\:characterString = "Auxiliary CTM AUX_CTMCH4 model input data" ;
                } // group gmd\:title

              group: gmd\:alternateTitle\#1 {

                // group attributes:
                		:gmx\:FileName = "S5P_OPER_AUX_CTMCH4_20240408T000000_20240409T000000_20231019T120000.nc" ;
                } // group gmd\:alternateTitle\#1

              group: gmd\:alternateTitle\#2 {

                // group attributes:
                		:gmx\:FileName = "S5P_OPER_AUX_CTMCH4_20240407T000000_20240408T000000_20231019T120000.nc" ;
                } // group gmd\:alternateTitle\#2
              } // group gmd\:sourceCitation
            } // group gmd\:source\#1

          group: gmd\:source\#2 {

            // group attributes:
            		:objectType = "gmi:LE_Source" ;
            		:gmd\:description = "Auxiliary CTM AUX_CTM_CO model input data" ;

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "N/A" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2024-04-09T12:47:23Z" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:title {

                // group attributes:
                		:gco\:characterString = "Auxiliary CTM AUX_CTM_CO model input data" ;
                } // group gmd\:title

              group: gmd\:alternateTitle\#1 {

                // group attributes:
                		:gmx\:FileName = "S5P_OPER_AUX_CTM_CO_20240101T000000_20250101T000000_20231019T120000.nc" ;
                } // group gmd\:alternateTitle\#1
              } // group gmd\:sourceCitation
            } // group gmd\:source\#2

          group: gmd\:source\#3 {

            // group attributes:
            		:objectType = "gmi:LE_Source" ;
            		:gmd\:description = "Auxiliary AUX_ISRF__ reference data" ;

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "N/A" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2024-04-09T12:47:23Z" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:title {

                // group attributes:
                		:gco\:characterString = "Auxiliary AUX_ISRF__ reference data" ;
                } // group gmd\:title

              group: gmd\:alternateTitle\#1 {

                // group attributes:
                		:gmx\:FileName = "S5P_OPER_AUX_ISRF___00000000T000000_99999999T999999_20210107T103220.nc" ;
                } // group gmd\:alternateTitle\#1
              } // group gmd\:sourceCitation
            } // group gmd\:source\#3

          group: gmd\:source\#4 {

            // group attributes:
            		:objectType = "gmi:LE_Source" ;
            		:gmd\:description = "Auxiliary ECMWF AUX_MET_2D Meteorological forecast data" ;

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "L4" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2024-04-09T12:47:23Z" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:title {

                // group attributes:
                		:gco\:characterString = "Auxiliary ECMWF AUX_MET_2D Meteorological forecast data" ;
                } // group gmd\:title

              group: gmd\:alternateTitle\#1 {

                // group attributes:
                		:gmx\:FileName = "S5P_OFFL_AUX_MET_2D_20240407T030000_20240407T120000_20240407T000000.nc" ;
                } // group gmd\:alternateTitle\#1

              group: gmd\:alternateTitle\#2 {

                // group attributes:
                		:gmx\:FileName = "S5P_OFFL_AUX_MET_2D_20240407T150000_20240408T000000_20240407T120000.nc" ;
                } // group gmd\:alternateTitle\#2
              } // group gmd\:sourceCitation
            } // group gmd\:source\#4

          group: gmd\:source\#5 {

            // group attributes:
            		:objectType = "gmi:LE_Source" ;
            		:gmd\:description = "Auxiliary ECMWF AUX_MET_QP Meteorological forecast data" ;

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "L4" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2024-04-09T12:47:23Z" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:title {

                // group attributes:
                		:gco\:characterString = "Auxiliary ECMWF AUX_MET_QP Meteorological forecast data" ;
                } // group gmd\:title

              group: gmd\:alternateTitle\#1 {

                // group attributes:
                		:gmx\:FileName = "S5P_OFFL_AUX_MET_QP_20240407T030000_20240407T120000_20240407T000000.nc" ;
                } // group gmd\:alternateTitle\#1

              group: gmd\:alternateTitle\#2 {

                // group attributes:
                		:gmx\:FileName = "S5P_OFFL_AUX_MET_QP_20240407T150000_20240408T000000_20240407T120000.nc" ;
                } // group gmd\:alternateTitle\#2
              } // group gmd\:sourceCitation
            } // group gmd\:source\#5

          group: gmd\:source\#6 {

            // group attributes:
            		:objectType = "gmi:LE_Source" ;
            		:gmd\:description = "Auxiliary ECMWF AUX_MET_TP Meteorological forecast data" ;

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "L4" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2024-04-09T12:47:23Z" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:title {

                // group attributes:
                		:gco\:characterString = "Auxiliary ECMWF AUX_MET_TP Meteorological forecast data" ;
                } // group gmd\:title

              group: gmd\:alternateTitle\#1 {

                // group attributes:
                		:gmx\:FileName = "S5P_OFFL_AUX_MET_TP_20240407T030000_20240407T120000_20240407T000000.nc" ;
                } // group gmd\:alternateTitle\#1

              group: gmd\:alternateTitle\#2 {

                // group attributes:
                		:gmx\:FileName = "S5P_OFFL_AUX_MET_TP_20240407T150000_20240408T000000_20240407T120000.nc" ;
                } // group gmd\:alternateTitle\#2
              } // group gmd\:sourceCitation
            } // group gmd\:source\#6

          group: gmd\:source\#7 {

            // group attributes:
            		:objectType = "gmi:LE_Source" ;
            		:gmd\:description = "Processor CFG_CH4__F configuration file" ;

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "N/A" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2024-04-09T12:47:23Z" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:title {

                // group attributes:
                		:gco\:characterString = "Processor CFG_CH4__F configuration file" ;
                } // group gmd\:title

              group: gmd\:alternateTitle\#1 {

                // group attributes:
                		:gmx\:FileName = "S5P_OPER_CFG_CH4__F_00000000T000000_99999999T999999_20230901T000000.cfg" ;
                } // group gmd\:alternateTitle\#1
              } // group gmd\:sourceCitation
            } // group gmd\:source\#7

          group: gmd\:source\#8 {

            // group attributes:
            		:objectType = "gmi:LE_Source" ;
            		:gmd\:description = "Processor CFG_CH4___ configuration file" ;

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "N/A" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2024-04-09T12:47:23Z" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:title {

                // group attributes:
                		:gco\:characterString = "Processor CFG_CH4___ configuration file" ;
                } // group gmd\:title

              group: gmd\:alternateTitle\#1 {

                // group attributes:
                		:gmx\:FileName = "S5P_OPER_CFG_CH4____00000000T000000_99999999T999999_20230901T000000.cfg" ;
                } // group gmd\:alternateTitle\#1
              } // group gmd\:sourceCitation
            } // group gmd\:source\#8

          group: gmd\:source\#9 {

            // group attributes:
            		:objectType = "gmi:LE_Source" ;
            		:gmd\:description = "TROPOMI L1B L1B_IR_SIR irradiance product" ;

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "L1B" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2024-04-09T12:47:23Z" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:title {

                // group attributes:
                		:gco\:characterString = "TROPOMI L1B L1B_IR_SIR irradiance product" ;
                } // group gmd\:title

              group: gmd\:alternateTitle\#1 {

                // group attributes:
                		:gmx\:FileName = "S5P_OFFL_L1B_IR_SIR_20240407T123946_20240407T142117_33598_03_020100_20240407T161058.nc" ;
                } // group gmd\:alternateTitle\#1
              } // group gmd\:sourceCitation
            } // group gmd\:source\#9

          group: gmd\:source\#10 {

            // group attributes:
            		:objectType = "gmi:LE_Source" ;
            		:gmd\:description = "TROPOMI L1B L1B_IR_UVN irradiance product" ;

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "L1B" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2024-04-09T12:47:23Z" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:title {

                // group attributes:
                		:gco\:characterString = "TROPOMI L1B L1B_IR_UVN irradiance product" ;
                } // group gmd\:title

              group: gmd\:alternateTitle\#1 {

                // group attributes:
                		:gmx\:FileName = "S5P_OFFL_L1B_IR_UVN_20240407T123946_20240407T142117_33598_03_020100_20240407T161058.nc" ;
                } // group gmd\:alternateTitle\#1
              } // group gmd\:sourceCitation
            } // group gmd\:source\#10

          group: gmd\:source\#11 {

            // group attributes:
            		:objectType = "gmi:LE_Source" ;
            		:gmd\:description = "TROPOMI L1B L1B_RA_BD6 radiance product" ;

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "L1B" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2024-04-09T12:47:23Z" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:title {

                // group attributes:
                		:gco\:characterString = "TROPOMI L1B L1B_RA_BD6 radiance product" ;
                } // group gmd\:title

              group: gmd\:alternateTitle\#1 {

                // group attributes:
                		:gmx\:FileName = "S5P_OFFL_L1B_RA_BD6_20240407T123946_20240407T142117_33598_03_020100_20240407T161058.nc" ;
                } // group gmd\:alternateTitle\#1
              } // group gmd\:sourceCitation
            } // group gmd\:source\#11

          group: gmd\:source\#12 {

            // group attributes:
            		:objectType = "gmi:LE_Source" ;
            		:gmd\:description = "TROPOMI L1B L1B_RA_BD7 radiance product" ;

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "L1B" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2024-04-09T12:47:23Z" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:title {

                // group attributes:
                		:gco\:characterString = "TROPOMI L1B L1B_RA_BD7 radiance product" ;
                } // group gmd\:title

              group: gmd\:alternateTitle\#1 {

                // group attributes:
                		:gmx\:FileName = "S5P_OFFL_L1B_RA_BD7_20240407T123946_20240407T142117_33598_03_020100_20240407T161058.nc" ;
                } // group gmd\:alternateTitle\#1
              } // group gmd\:sourceCitation
            } // group gmd\:source\#12

          group: gmd\:source\#13 {

            // group attributes:
            		:objectType = "gmi:LE_Source" ;
            		:gmd\:description = "TROPOMI L1B L1B_RA_BD8 radiance product" ;

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "L1B" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2024-04-09T12:47:23Z" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:title {

                // group attributes:
                		:gco\:characterString = "TROPOMI L1B L1B_RA_BD8 radiance product" ;
                } // group gmd\:title

              group: gmd\:alternateTitle\#1 {

                // group attributes:
                		:gmx\:FileName = "S5P_OFFL_L1B_RA_BD8_20240407T123946_20240407T142117_33598_03_020100_20240407T161058.nc" ;
                } // group gmd\:alternateTitle\#1
              } // group gmd\:sourceCitation
            } // group gmd\:source\#13

          group: gmd\:source\#14 {

            // group attributes:
            		:objectType = "gmi:LE_Source" ;
            		:gmd\:description = "TROPOMI L2 L2__CH4CLD product" ;

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "N/A" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2024-04-09T12:47:23Z" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:title {

                // group attributes:
                		:gco\:characterString = "TROPOMI L2 L2__CH4CLD product" ;
                } // group gmd\:title

              group: gmd\:alternateTitle\#1 {

                // group attributes:
                		:gmx\:FileName = "S5P_OFFL_L2__CH4CLD_20240407T123946_20240407T142117_33598_03_020600_20240409T045645.nc" ;
                } // group gmd\:alternateTitle\#1
              } // group gmd\:sourceCitation
            } // group gmd\:source\#14

          group: gmd\:source\#15 {

            // group attributes:
            		:objectType = "gmi:LE_Source" ;
            		:gmd\:description = "TROPOMI L2 L2__CO____ product" ;

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "N/A" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2024-04-09T12:47:23Z" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:title {

                // group attributes:
                		:gco\:characterString = "TROPOMI L2 L2__CO____ product" ;
                } // group gmd\:title

              group: gmd\:alternateTitle\#1 {

                // group attributes:
                		:gmx\:FileName = "S5P_OFFL_L2__CO_____20240407T123946_20240407T142117_33598_03_020600_20240409T023051.nc" ;
                } // group gmd\:alternateTitle\#1
              } // group gmd\:sourceCitation
            } // group gmd\:source\#15

          group: gmd\:source\#16 {

            // group attributes:
            		:objectType = "gmi:LE_Source" ;
            		:gmd\:description = "TROPOMI L2 L2__FRESCO product" ;

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "N/A" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2024-04-09T12:47:23Z" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:title {

                // group attributes:
                		:gco\:characterString = "TROPOMI L2 L2__FRESCO product" ;
                } // group gmd\:title

              group: gmd\:alternateTitle\#1 {

                // group attributes:
                		:gmx\:FileName = "S5P_OFFL_L2__FRESCO_20240407T123946_20240407T142117_33598_03_020600_20240409T023052.nc" ;
                } // group gmd\:alternateTitle\#1
              } // group gmd\:sourceCitation
            } // group gmd\:source\#16

          group: gmd\:source\#17 {

            // group attributes:
            		:objectType = "gmi:LE_Source" ;
            		:gmd\:description = "TROPOMI L2 L2__NP_BD6 product" ;

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "N/A" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2024-04-09T12:47:23Z" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:title {

                // group attributes:
                		:gco\:characterString = "TROPOMI L2 L2__NP_BD6 product" ;
                } // group gmd\:title

              group: gmd\:alternateTitle\#1 {

                // group attributes:
                		:gmx\:FileName = "S5P_OFFL_L2__NP_BD6_20240407T123946_20240407T142117_33598_03_020000_20240409T023051.nc" ;
                } // group gmd\:alternateTitle\#1
              } // group gmd\:sourceCitation
            } // group gmd\:source\#17

          group: gmd\:source\#18 {

            // group attributes:
            		:objectType = "gmi:LE_Source" ;
            		:gmd\:description = "TROPOMI L2 L2__NP_BD7 product" ;

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "N/A" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2024-04-09T12:47:23Z" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:title {

                // group attributes:
                		:gco\:characterString = "TROPOMI L2 L2__NP_BD7 product" ;
                } // group gmd\:title

              group: gmd\:alternateTitle\#1 {

                // group attributes:
                		:gmx\:FileName = "S5P_OFFL_L2__NP_BD7_20240407T123946_20240407T142117_33598_03_020000_20240409T023051.nc" ;
                } // group gmd\:alternateTitle\#1
              } // group gmd\:sourceCitation
            } // group gmd\:source\#18

          group: gmd\:source\#19 {

            // group attributes:
            		:objectType = "gmi:LE_Source" ;
            		:gmd\:description = "Auxiliary LUT_CH4AER algorithm lookup table" ;

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "N/A" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2024-04-09T12:47:23Z" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:title {

                // group attributes:
                		:gco\:characterString = "Auxiliary LUT_CH4AER algorithm lookup table" ;
                } // group gmd\:title

              group: gmd\:alternateTitle\#1 {

                // group attributes:
                		:gmx\:FileName = "S5P_OPER_LUT_CH4AER_00000000T000000_99999999T999999_20151008T180555.nc" ;
                } // group gmd\:alternateTitle\#1
              } // group gmd\:sourceCitation
            } // group gmd\:source\#19

          group: gmd\:source\#20 {

            // group attributes:
            		:objectType = "gmi:LE_Source" ;
            		:gmd\:description = "Auxiliary LUT_CH4CIR algorithm lookup table" ;

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "N/A" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2024-04-09T12:47:23Z" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:title {

                // group attributes:
                		:gco\:characterString = "Auxiliary LUT_CH4CIR algorithm lookup table" ;
                } // group gmd\:title

              group: gmd\:alternateTitle\#1 {

                // group attributes:
                		:gmx\:FileName = "S5P_OPER_LUT_CH4CIR_00000000T000000_99999999T999999_20151016T113037.nc" ;
                } // group gmd\:alternateTitle\#1
              } // group gmd\:sourceCitation
            } // group gmd\:source\#20

          group: gmd\:source\#21 {

            // group attributes:
            		:objectType = "gmi:LE_Source" ;
            		:gmd\:description = "Auxiliary LUT_CH4RFC algorithm lookup table" ;

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "N/A" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2024-04-09T12:47:23Z" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:title {

                // group attributes:
                		:gco\:characterString = "Auxiliary LUT_CH4RFC algorithm lookup table" ;
                } // group gmd\:title

              group: gmd\:alternateTitle\#1 {

                // group attributes:
                		:gmx\:FileName = "S5P_OPER_LUT_CH4RFC_00000000T000000_99999999T999999_20230720T134206.zip" ;
                } // group gmd\:alternateTitle\#1
              } // group gmd\:sourceCitation
            } // group gmd\:source\#21

          group: gmd\:source\#22 {

            // group attributes:
            		:objectType = "gmi:LE_Source" ;
            		:gmd\:description = "Auxiliary REF_DEM___ reference data" ;

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "N/A" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2024-04-09T12:47:23Z" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:title {

                // group attributes:
                		:gco\:characterString = "Auxiliary REF_DEM___ reference data" ;
                } // group gmd\:title

              group: gmd\:alternateTitle\#1 {

                // group attributes:
                		:gmx\:FileName = "S5P_OPER_REF_DEM____20190404T150000_99999999T999999_20190405T143622.nc" ;
                } // group gmd\:alternateTitle\#1
              } // group gmd\:sourceCitation
            } // group gmd\:source\#22

          group: gmd\:source\#23 {

            // group attributes:
            		:objectType = "gmi:LE_Source" ;
            		:gmd\:description = "Auxiliary REF_SOLAR_ reference data" ;

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "N/A" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2024-04-09T12:47:23Z" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:title {

                // group attributes:
                		:gco\:characterString = "Auxiliary REF_SOLAR_ reference data" ;
                } // group gmd\:title

              group: gmd\:alternateTitle\#1 {

                // group attributes:
                		:gmx\:FileName = "S5P_OPER_REF_SOLAR__00000000T000000_99999999T999999_20210107T132455.nc" ;
                } // group gmd\:alternateTitle\#1
              } // group gmd\:sourceCitation
            } // group gmd\:source\#23

          group: gmd\:source\#24 {

            // group attributes:
            		:objectType = "gmi:LE_Source" ;
            		:gmd\:description = "Auxiliary REF_XS_CH4 reference data" ;

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "N/A" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2024-04-09T12:47:23Z" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:title {

                // group attributes:
                		:gco\:characterString = "Auxiliary REF_XS_CH4 reference data" ;
                } // group gmd\:title

              group: gmd\:alternateTitle\#1 {

                // group attributes:
                		:gmx\:FileName = "S5P_OPER_REF_XS_CH4_00000000T000000_99999999T999999_20200710T082601.nc" ;
                } // group gmd\:alternateTitle\#1
              } // group gmd\:sourceCitation
            } // group gmd\:source\#24
          } // group gmd\:processStep
        } // group gmd\:lineage
      } // group gmd\:dataQualityInfo

    group: gmi\:acquisitionInformation {

      // group attributes:
      		:objectType = "gmi:MI_AcquisitionInformation" ;

      group: gmi\:platform {

        // group attributes:
        		:gmi\:description = "Sentinel 5 Precursor" ;
        		:objectType = "gmi:MI_Platform" ;

        group: gmi\:identifier {

          // group attributes:
          		:gmd\:code = "S5P" ;
          		:gmd\:codeSpace = "http://www.esa.int/" ;
          		:objectType = "gmd:RS_Identifier" ;
          } // group gmi\:identifier

        group: gmi\:instrument {

          // group attributes:
          		:objectType = "gmi:MI_Instrument" ;
          		:gmi\:type = "UV-VIS-NIR-SWIR imaging spectrometer" ;

          group: gmi\:identifier {

            // group attributes:
            		:gmd\:code = "TROPOMI" ;
            		:gmd\:codeSpace = "http://www.esa.int/" ;
            		:objectType = "gmd:RS_Identifier" ;
            } // group gmi\:identifier
          } // group gmi\:instrument
        } // group gmi\:platform
      } // group gmi\:acquisitionInformation
    } // group ISO_METADATA

  group: EOP_METADATA {

    // group attributes:
    		:gml\:id = "S5P_OFFL_L2__CH4____20240407T123946_20240407T142117_33598_03_020600_20240409T045638.ID" ;
    		:objectType = "atm:EarthObservation" ;

    group: om\:phenomenonTime {

      // group attributes:
      		:gml\:beginPosition = "2024-04-07T13:01:21Z" ;
      		:gml\:endPosition = "2024-04-07T13:53:37Z" ;
      		:objectType = "gml:TimePeriod" ;
      } // group om\:phenomenonTime

    group: om\:procedure {

      // group attributes:
      		:gml\:id = "S5P_OFFL_L2__CH4____20240407T123946_20240407T142117_33598_03_020600_20240409T045638.EOE" ;
      		:objectType = "eop:EarthObservationEquipment" ;

      group: eop\:platform {

        // group attributes:
        		:eop\:shortName = "Sentinel-5p" ;
        		:objectType = "eop:Platform" ;
        } // group eop\:platform

      group: eop\:instrument {

        // group attributes:
        		:eop\:shortName = "TROPOMI" ;
        		:objectType = "eop:Instrument" ;
        } // group eop\:instrument

      group: eop\:sensor {

        // group attributes:
        		:eop\:sensorType = "ATMOSPHERIC" ;
        		:objectType = "eop:Sensor" ;
        } // group eop\:sensor

      group: eop\:acquisitionParameters {

        // group attributes:
        		:eop\:orbitNumber = 33598 ;
        		:objectType = "eop:Acquisition" ;
        } // group eop\:acquisitionParameters
      } // group om\:procedure

    group: om\:observedProperty {

      // group attributes:
      		:nilReason = "inapplicable" ;
      } // group om\:observedProperty

    group: om\:featureOfInterest {

      // group attributes:
      		:objectType = "eop:FootPrint" ;
      		:gml\:id = "S5P_OFFL_L2__CH4____20240407T123946_20240407T142117_33598_03_020600_20240409T045638.FP" ;

      group: eop\:multiExtentOf {

        // group attributes:
        		:objectType = "gml:MultiSurface" ;

        group: gml\:surfaceMembers {

          // group attributes:
          		:objectType = "gml:Polygon" ;

          group: gml\:exterior {

            // group attributes:
            		:gml\:posList = "69.12326 -96.52095 68.9921 -94.0861 68.86768 -91.2714 68.70395 -87.12199 68.43766 -83.05291 68.07201 -79.09739 67.61219 -75.283356 67.06428 -71.63077 66.433426 -68.155045 65.727 -64.863235 64.95094 -61.758682 64.11166 -58.839714 63.21494 -56.10169 62.26636 -53.53706 61.271183 -51.137142 60.234016 -48.892162 59.15911 -46.791767 58.05016 -44.826317 56.910427 -42.98577 55.743427 -41.260048 54.551414 -39.64084 53.336998 -38.11939 52.10234 -36.687958 50.84924 -35.33934 49.57952 -34.06696 48.294548 -32.864838 46.995846 -31.727276 45.68447 -30.649435 44.361584 -29.62661 43.028168 -28.65449 41.68505 -27.729483 40.332916 -26.848196 38.972782 -26.007145 37.60501 -25.203585 36.230232 -24.43517 34.84901 -23.699062 33.46196 -22.9933 32.069298 -22.31575 30.671553 -21.664774 29.269096 -21.038534 27.86219 -20.43558 26.451256 -19.854311 25.036455 -19.2936 23.618092 -18.752457 22.196503 -18.229338 20.771818 -17.723442 19.344297 -17.234015 17.914246 -16.759632 16.481695 -16.300047 15.046912 -15.854254 13.610022 -15.42169 12.171148 -15.001694 10.7305565 -14.593701 9.288325 -14.197052 7.844606 -13.811342 6.399445 -13.436193 4.9529796 -13.071237 3.5054948 -12.715716 2.056944 -12.369523 0.60745215 -12.032404 -0.8428004 -11.703914 -2.2938066 -11.383875 -3.7453773 -11.071796 -5.197478 -10.767557 -6.6501603 -10.471336 -8.103019 -10.182347 -9.55626 -9.900891 -11.009554 -9.626229 -12.4630375 -9.358874 -13.916575 -9.098447 -15.370095 -8.844885 -16.82345 -8.598179 -18.276707 -8.358217 -19.72974 -8.124872 -21.182499 -7.8985233 -22.634861 -7.678618 -24.086777 -7.465518 -25.538235 -7.2592893 -26.989267 -7.059948 -28.439674 -6.8678403 -29.889502 -6.682653 -31.338615 -6.505009 -32.787018 -6.334882 -34.23472 -6.1726823 -35.681602 -6.018626 -37.127575 -5.8727093 -38.572773 -5.7362585 -40.01691 -5.6086483 -41.460114 -5.4909673 -42.902348 -5.383861 -44.34349 -5.287823 -45.78353 -5.2034283 -47.22245 -5.13245 -48.660156 -5.0750704 -50.096634 -5.0329905 -51.531773 -5.007261 -52.96554 -4.999523 -54.39791 -5.0120163 -55.828766 -5.046724 -57.258034 -5.1065807 -58.685528 -5.1945086 -60.111244 -5.3141966 -61.53498 -5.4701643 -62.95653 -5.6681566 -64.37574 -5.914327 -65.792274 -6.2169905 -67.205765 -6.585456 -68.61589 -7.0346236 -70.021996 -7.5789742 -71.42331 -8.239928 -72.81896 -9.046077 -74.20753 -10.034298 -75.58711 -11.255124 -76.955185 -12.779777 -78.30788 -14.711452 -79.63933 -17.20201 -80.940346 -20.48162 -82.196175 -24.908434 -83.381 -31.055166 -84.44982 -39.801342 -85.32229 -52.322144 -85.872116 -69.35114 -85.96579 -89.23881 -85.57413 -107.71778 -84.80586 -121.915825 -84.32533 -127.37689 -84.61155 -129.5894 -86.26667 -154.16481 -86.62555 168.91461 -86.17712 149.70721 -85.32004 135.04347 -84.65357 128.58513 -83.79734 123.021065 -83.18459 120.16023 -82.39927 117.37243 -81.825935 115.786194 -81.06929 114.117584 -80.49823 113.10717 -79.71702 111.99399 -79.1045 111.29605 -78.23123 110.51073 -77.51515 110.013824 -76.44068 109.457565 -75.50644 109.11234 -73.99777 108.73895 -72.55751 108.517204 -69.87725 108.28098 -68.63999 108.20952 -68.86911 104.10728 -68.99504 99.93759 -69.01601 95.73987 -68.931725 91.5541 -68.743126 87.42037 -68.453316 83.375206 -68.06614 79.450485 -67.58648 75.67274 -67.02021 72.060585 -66.37354 68.62667 -65.65293 65.37805 -64.864655 62.316147 -64.014786 59.438873 -63.1092 56.740433 -62.1532 54.213306 -61.151844 51.848297 -60.109577 49.63584 -59.030815 47.565193 -57.91874 45.62712 -56.77701 43.811134 -55.60827 42.108334 -54.415405 40.509342 -53.20077 39.006058 -51.96629 37.59109 -50.71379 36.257175 -49.44485 34.998173 -48.161076 33.80803 -46.86386 32.6809 -45.554195 31.612541 -44.233177 30.597982 -42.90178 29.633245 -41.560883 28.7145 -40.211098 27.838762 -38.85333 27.002571 -37.488033 26.203236 -36.11591 25.43806 -34.737293 24.704924 -33.35287 24.001442 -31.962915 23.325813 -30.567896 22.6761 -29.168053 22.050915 -27.763897 21.448427 -26.355658 20.86747 -24.943605 20.30639 -23.527925 19.764442 -22.109062 19.240267 -20.68719 18.733051 -19.26225 18.24198 -17.834806 17.765865 -16.404867 17.30402 -14.972613 16.855686 -13.5382595 16.420498 -12.101926 15.997358 -10.663737 15.586139 -9.223851 15.1859455 -7.782439 14.796269 -6.3396125 14.417082 -4.895427 14.047611 -3.450113 13.687472 -2.0036685 13.336456 -0.5562642 12.994084 0.89207447 12.660093 2.3410919 12.333932 3.7909138 12.015948 5.2413144 11.705307 6.692206 11.402052 8.143573 11.105971 9.595263 10.816896 11.047319 10.534819 12.499652 10.259289 13.952056 9.990306 15.404554 9.727688 16.857092 9.471441 18.309643 9.221598 19.762098 8.977995 21.214369 8.740265 22.666468 8.509207 24.118393 8.284123 25.569899 8.065376 27.021118 7.852739 28.472 7.646652 29.92251 7.4465227 31.372461 7.2536473 32.821968 7.0672526 34.270992 6.887798 35.719368 6.7155194 37.16717 6.550701 38.614338 6.393722 40.06086 6.2448573 41.506695 6.1044188 42.951824 5.972929 44.396248 5.8515277 45.83986 5.739734 47.282642 5.639565 48.7246 5.551 50.16572 5.4754996 51.60594 5.4140086 53.04517 5.368121 54.4834 5.3393207 55.920586 5.329705 57.356674 5.341325 58.7916 5.3769507 60.225357 5.439257 61.657753 5.532945 63.088596 5.6622677 64.51782 5.8330317 65.94532 6.0518312 67.37069 6.328257 68.79367 6.6737347 70.21398 7.1015344 71.630875 7.63117 73.04383 8.28766 74.45169 9.104776 75.85312 10.130339 77.24618 11.428328 78.627846 13.099217 79.99347 15.290404 81.33562 18.238403 82.64159 22.326872 83.88807 28.224384 85.03025 37.082226 85.978584 50.74104 86.5691 71.113495 86.188515 110.07581 85.7742 119.710754 86.01269 122.72938 87.19441 157.42668 86.85943 -160.9204 86.13021 -144.85469 85.126816 -133.49129 84.42676 -128.35394 83.56847 -123.62431 82.970314 -120.9771 82.21566 -118.1496 81.67048 -116.37208 80.95599 -114.29774 80.41942 -112.89214 79.68786 -111.143585 79.115585 -109.887115 78.30068 -108.236496 77.632515 -106.98647 76.62838 -105.2584 75.75219 -103.88214 74.32772 -101.87871 72.953415 -100.191795 70.34922 -97.55307 69.12326 -96.52095 69.12326 -96.52095" ;
            		:objectType = "gml:LinearRing" ;
            } // group gml\:exterior
          } // group gml\:surfaceMembers
        } // group eop\:multiExtentOf
      } // group om\:featureOfInterest

    group: eop\:metaDataProperty {

      // group attributes:
      		:objectType = "eop:EarthObservationMetaData" ;
      		:eop\:acquisitionType = "NOMINAL" ;
      		:eop\:identifier = "S5P_OFFL_L2__CH4____20240407T123946_20240407T142117_33598_03_020600_20240409T045638" ;
      		:eop\:doi = "10.5270/S5P-3lcdqiv" ;
      		:eop\:parentIdentifier = "urn:ogc:def:EOP:ESA:SENTINEL.S5P_TROP_L2__CH4___" ;
      		:eop\:productType = "S5P_OFFL_CH4___" ;
      		:eop\:status = "ACQUIRED" ;
      		:eop\:productQualityStatus = "NOMINAL" ;
      		:eop\:productQualityDegradationTag = "NOT APPLICABLE" ;

      group: eop\:processing {

        // group attributes:
        		:objectType = "eop:ProcessingInformation" ;
        		:eop\:processingCenter = "PDGS-OP" ;
        		:eop\:processingDate = "2024-04-09" ;
        		:eop\:processingLevel = "L2" ;
        		:eop\:processorName = "TROPNLL2DP" ;
        		:eop\:processorVersion = "2.6.0" ;
        		:eop\:nativeProductFormat = "netCDF-4" ;
        		:eop\:processingMode = "OFFL" ;
        } // group eop\:processing
      } // group eop\:metaDataProperty
    } // group EOP_METADATA

  group: ESA_METADATA {

    group: earth_explorer_header {

      // group attributes:
      		:objectType = "Earth_Explorer_Header" ;

      group: fixed_header {

        // group attributes:
        		:objectType = "Fixed_Header" ;
        		:File_Name = "S5P_OFFL_L2__CH4____20240407T123946_20240407T142117_33598_03_020600_20240409T045638" ;
        		:File_Description = "Dry-air mixing ratio of methane for cloud-free observations with a spatial resolution of 5.5x7.0 km2 observed at about 13:30 local solar time from spectra measured by TROPOMI" ;
        		:Notes = "" ;
        		:Mission = "S5P" ;
        		:File_Class = "OFFL" ;
        		:File_Type = "L2__CH4___" ;
        		:File_Version = 1 ;

        group: validity_period {

          // group attributes:
          		:objectType = "Validity_Period" ;
          		:Validity_Start = "UTC=2024-04-07T13:01:21" ;
          		:Validity_Stop = "UTC=2024-04-07T13:53:37" ;
          } // group validity_period

        group: source {

          // group attributes:
          		:objectType = "Source" ;
          		:System = "PDGS-OP" ;
          		:Creator = "TROPNLL2DP" ;
          		:Creator_Version = "2.6.0" ;
          		:Creation_Date = "UTC=2024-04-09T05:04:45" ;
          } // group source
        } // group fixed_header

      group: variable_header {

        // group attributes:
        		:objectType = "Variable_Header" ;

        group: gmd\:lineage {

          // group attributes:
          		:objectType = "gmd:LI_Lineage" ;
          		:gmd\:statement = "L2 CH4___ dataset produced by PDGS-OP from the S5P/TROPOMI L1B product" ;

          group: gmd\:processStep {

            // group attributes:
            		:objectType = "gmi:LE_ProcessStep" ;
            		:gmd\:description = "Processing of L1b to L2 CH4___ data for orbit 33598 using the KNMI/SRON processor version 2.6.0" ;

            group: gmi\:output {

              // group attributes:
              		:gmd\:description = "TROPOMI/S5P Methane 1-Orbit L2 Swath 5.5x7.0km" ;
              		:objectType = "gmi:LE_Source" ;

              group: gmd\:sourceCitation {

                // group attributes:
                		:gmd\:title = "S5P_OFFL_L2__CH4____20240407T123946_20240407T142117_33598_03_020600_20240409T045638" ;
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2024-04-09" ;
                  		:objectType = "gmd:CI_DateTime" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:identifier {

                  // group attributes:
                  		:gmd\:code = "L2__CH4___" ;
                  		:objectType = "gmd:MD_Identifier" ;
                  } // group gmd\:identifier
                } // group gmd\:sourceCitation

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "L2" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel
              } // group gmi\:output

            group: gmi\:processingInformation {

              // group attributes:
              		:objectType = "gmi:LE_Processing" ;

              group: gmi\:identifier {

                // group attributes:
                		:gmd\:code = "KNMI/SRON L2 CH4___ processor, version 2.6.0" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:identifier

              group: gmi\:softwareReference {

                // group attributes:
                		:gmd\:title = "TROPNLL2DP processor" ;
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2023-09-28T07:04:00Z" ;
                  		:objectType = "gmd:CI_DateTime" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date
                } // group gmi\:softwareReference

              group: gmi\:documentation\#1 {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;
                		:gmd\:title = "Algorithm Theoretical Baseline Document for Sentinel-5 Precursor Methane Retrieval; SRON-S5P-LEV2-RP-001; release 1.0" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2015-11-30" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "revision" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date
                } // group gmi\:documentation\#1

              group: gmi\:documentation\#2 {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;
                		:gmd\:title = "Sentinel-5 precursor/TROPOMI Level 2 Product User Manual Methane; SRON-S5P-LEV2-MA-001; release 1.0" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2015-11-30" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "revision" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date
                } // group gmi\:documentation\#2
              } // group gmi\:processingInformation

            group: gmi\:report {

              // group attributes:
              		:gmi\:description = "Sentinel 5-precursor TROPOMI L1b processed to L2 data using the KNMI/SRON L2 CH4___ processor" ;
              		:gmi\:fileType = "netCDF-4" ;
              		:gmi\:name = "S5P_OFFL_L2__CH4____20240407T123946_20240407T142117_33598_03_020600_20240409T045638.nc" ;
              		:objectType = "gmi:LE_ProcessStepReport" ;
              } // group gmi\:report

            group: gmd\:source\#1 {

              // group attributes:
              		:objectType = "gmi:LE_Source" ;
              		:gmd\:description = "Auxiliary CTM AUX_CTMCH4 model input data" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "N/A" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2024-04-09T12:47:23Z" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "Auxiliary CTM AUX_CTMCH4 model input data" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_OPER_AUX_CTMCH4_20240408T000000_20240409T000000_20231019T120000.nc" ;
                  } // group gmd\:alternateTitle\#1

                group: gmd\:alternateTitle\#2 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_OPER_AUX_CTMCH4_20240407T000000_20240408T000000_20231019T120000.nc" ;
                  } // group gmd\:alternateTitle\#2
                } // group gmd\:sourceCitation
              } // group gmd\:source\#1

            group: gmd\:source\#2 {

              // group attributes:
              		:objectType = "gmi:LE_Source" ;
              		:gmd\:description = "Auxiliary CTM AUX_CTM_CO model input data" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "N/A" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2024-04-09T12:47:23Z" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "Auxiliary CTM AUX_CTM_CO model input data" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_OPER_AUX_CTM_CO_20240101T000000_20250101T000000_20231019T120000.nc" ;
                  } // group gmd\:alternateTitle\#1
                } // group gmd\:sourceCitation
              } // group gmd\:source\#2

            group: gmd\:source\#3 {

              // group attributes:
              		:objectType = "gmi:LE_Source" ;
              		:gmd\:description = "Auxiliary AUX_ISRF__ reference data" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "N/A" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2024-04-09T12:47:23Z" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "Auxiliary AUX_ISRF__ reference data" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_OPER_AUX_ISRF___00000000T000000_99999999T999999_20210107T103220.nc" ;
                  } // group gmd\:alternateTitle\#1
                } // group gmd\:sourceCitation
              } // group gmd\:source\#3

            group: gmd\:source\#4 {

              // group attributes:
              		:objectType = "gmi:LE_Source" ;
              		:gmd\:description = "Auxiliary ECMWF AUX_MET_2D Meteorological forecast data" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "L4" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2024-04-09T12:47:23Z" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "Auxiliary ECMWF AUX_MET_2D Meteorological forecast data" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_OFFL_AUX_MET_2D_20240407T030000_20240407T120000_20240407T000000.nc" ;
                  } // group gmd\:alternateTitle\#1

                group: gmd\:alternateTitle\#2 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_OFFL_AUX_MET_2D_20240407T150000_20240408T000000_20240407T120000.nc" ;
                  } // group gmd\:alternateTitle\#2
                } // group gmd\:sourceCitation
              } // group gmd\:source\#4

            group: gmd\:source\#5 {

              // group attributes:
              		:objectType = "gmi:LE_Source" ;
              		:gmd\:description = "Auxiliary ECMWF AUX_MET_QP Meteorological forecast data" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "L4" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2024-04-09T12:47:23Z" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "Auxiliary ECMWF AUX_MET_QP Meteorological forecast data" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_OFFL_AUX_MET_QP_20240407T030000_20240407T120000_20240407T000000.nc" ;
                  } // group gmd\:alternateTitle\#1

                group: gmd\:alternateTitle\#2 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_OFFL_AUX_MET_QP_20240407T150000_20240408T000000_20240407T120000.nc" ;
                  } // group gmd\:alternateTitle\#2
                } // group gmd\:sourceCitation
              } // group gmd\:source\#5

            group: gmd\:source\#6 {

              // group attributes:
              		:objectType = "gmi:LE_Source" ;
              		:gmd\:description = "Auxiliary ECMWF AUX_MET_TP Meteorological forecast data" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "L4" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2024-04-09T12:47:23Z" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "Auxiliary ECMWF AUX_MET_TP Meteorological forecast data" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_OFFL_AUX_MET_TP_20240407T030000_20240407T120000_20240407T000000.nc" ;
                  } // group gmd\:alternateTitle\#1

                group: gmd\:alternateTitle\#2 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_OFFL_AUX_MET_TP_20240407T150000_20240408T000000_20240407T120000.nc" ;
                  } // group gmd\:alternateTitle\#2
                } // group gmd\:sourceCitation
              } // group gmd\:source\#6

            group: gmd\:source\#7 {

              // group attributes:
              		:objectType = "gmi:LE_Source" ;
              		:gmd\:description = "Processor CFG_CH4__F configuration file" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "N/A" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2024-04-09T12:47:23Z" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "Processor CFG_CH4__F configuration file" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_OPER_CFG_CH4__F_00000000T000000_99999999T999999_20230901T000000.cfg" ;
                  } // group gmd\:alternateTitle\#1
                } // group gmd\:sourceCitation
              } // group gmd\:source\#7

            group: gmd\:source\#8 {

              // group attributes:
              		:objectType = "gmi:LE_Source" ;
              		:gmd\:description = "Processor CFG_CH4___ configuration file" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "N/A" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2024-04-09T12:47:23Z" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "Processor CFG_CH4___ configuration file" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_OPER_CFG_CH4____00000000T000000_99999999T999999_20230901T000000.cfg" ;
                  } // group gmd\:alternateTitle\#1
                } // group gmd\:sourceCitation
              } // group gmd\:source\#8

            group: gmd\:source\#9 {

              // group attributes:
              		:objectType = "gmi:LE_Source" ;
              		:gmd\:description = "TROPOMI L1B L1B_IR_SIR irradiance product" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "L1B" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2024-04-09T12:47:23Z" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "TROPOMI L1B L1B_IR_SIR irradiance product" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_OFFL_L1B_IR_SIR_20240407T123946_20240407T142117_33598_03_020100_20240407T161058.nc" ;
                  } // group gmd\:alternateTitle\#1
                } // group gmd\:sourceCitation
              } // group gmd\:source\#9

            group: gmd\:source\#10 {

              // group attributes:
              		:objectType = "gmi:LE_Source" ;
              		:gmd\:description = "TROPOMI L1B L1B_IR_UVN irradiance product" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "L1B" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2024-04-09T12:47:23Z" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "TROPOMI L1B L1B_IR_UVN irradiance product" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_OFFL_L1B_IR_UVN_20240407T123946_20240407T142117_33598_03_020100_20240407T161058.nc" ;
                  } // group gmd\:alternateTitle\#1
                } // group gmd\:sourceCitation
              } // group gmd\:source\#10

            group: gmd\:source\#11 {

              // group attributes:
              		:objectType = "gmi:LE_Source" ;
              		:gmd\:description = "TROPOMI L1B L1B_RA_BD6 radiance product" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "L1B" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2024-04-09T12:47:23Z" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "TROPOMI L1B L1B_RA_BD6 radiance product" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_OFFL_L1B_RA_BD6_20240407T123946_20240407T142117_33598_03_020100_20240407T161058.nc" ;
                  } // group gmd\:alternateTitle\#1
                } // group gmd\:sourceCitation
              } // group gmd\:source\#11

            group: gmd\:source\#12 {

              // group attributes:
              		:objectType = "gmi:LE_Source" ;
              		:gmd\:description = "TROPOMI L1B L1B_RA_BD7 radiance product" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "L1B" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2024-04-09T12:47:23Z" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "TROPOMI L1B L1B_RA_BD7 radiance product" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_OFFL_L1B_RA_BD7_20240407T123946_20240407T142117_33598_03_020100_20240407T161058.nc" ;
                  } // group gmd\:alternateTitle\#1
                } // group gmd\:sourceCitation
              } // group gmd\:source\#12

            group: gmd\:source\#13 {

              // group attributes:
              		:objectType = "gmi:LE_Source" ;
              		:gmd\:description = "TROPOMI L1B L1B_RA_BD8 radiance product" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "L1B" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2024-04-09T12:47:23Z" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "TROPOMI L1B L1B_RA_BD8 radiance product" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_OFFL_L1B_RA_BD8_20240407T123946_20240407T142117_33598_03_020100_20240407T161058.nc" ;
                  } // group gmd\:alternateTitle\#1
                } // group gmd\:sourceCitation
              } // group gmd\:source\#13

            group: gmd\:source\#14 {

              // group attributes:
              		:objectType = "gmi:LE_Source" ;
              		:gmd\:description = "TROPOMI L2 L2__CH4CLD product" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "N/A" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2024-04-09T12:47:23Z" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "TROPOMI L2 L2__CH4CLD product" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_OFFL_L2__CH4CLD_20240407T123946_20240407T142117_33598_03_020600_20240409T045645.nc" ;
                  } // group gmd\:alternateTitle\#1
                } // group gmd\:sourceCitation
              } // group gmd\:source\#14

            group: gmd\:source\#15 {

              // group attributes:
              		:objectType = "gmi:LE_Source" ;
              		:gmd\:description = "TROPOMI L2 L2__CO____ product" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "N/A" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2024-04-09T12:47:23Z" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "TROPOMI L2 L2__CO____ product" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_OFFL_L2__CO_____20240407T123946_20240407T142117_33598_03_020600_20240409T023051.nc" ;
                  } // group gmd\:alternateTitle\#1
                } // group gmd\:sourceCitation
              } // group gmd\:source\#15

            group: gmd\:source\#16 {

              // group attributes:
              		:objectType = "gmi:LE_Source" ;
              		:gmd\:description = "TROPOMI L2 L2__FRESCO product" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "N/A" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2024-04-09T12:47:23Z" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "TROPOMI L2 L2__FRESCO product" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_OFFL_L2__FRESCO_20240407T123946_20240407T142117_33598_03_020600_20240409T023052.nc" ;
                  } // group gmd\:alternateTitle\#1
                } // group gmd\:sourceCitation
              } // group gmd\:source\#16

            group: gmd\:source\#17 {

              // group attributes:
              		:objectType = "gmi:LE_Source" ;
              		:gmd\:description = "TROPOMI L2 L2__NP_BD6 product" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "N/A" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2024-04-09T12:47:23Z" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "TROPOMI L2 L2__NP_BD6 product" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_OFFL_L2__NP_BD6_20240407T123946_20240407T142117_33598_03_020000_20240409T023051.nc" ;
                  } // group gmd\:alternateTitle\#1
                } // group gmd\:sourceCitation
              } // group gmd\:source\#17

            group: gmd\:source\#18 {

              // group attributes:
              		:objectType = "gmi:LE_Source" ;
              		:gmd\:description = "TROPOMI L2 L2__NP_BD7 product" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "N/A" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2024-04-09T12:47:23Z" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "TROPOMI L2 L2__NP_BD7 product" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_OFFL_L2__NP_BD7_20240407T123946_20240407T142117_33598_03_020000_20240409T023051.nc" ;
                  } // group gmd\:alternateTitle\#1
                } // group gmd\:sourceCitation
              } // group gmd\:source\#18

            group: gmd\:source\#19 {

              // group attributes:
              		:objectType = "gmi:LE_Source" ;
              		:gmd\:description = "Auxiliary LUT_CH4AER algorithm lookup table" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "N/A" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2024-04-09T12:47:23Z" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "Auxiliary LUT_CH4AER algorithm lookup table" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_OPER_LUT_CH4AER_00000000T000000_99999999T999999_20151008T180555.nc" ;
                  } // group gmd\:alternateTitle\#1
                } // group gmd\:sourceCitation
              } // group gmd\:source\#19

            group: gmd\:source\#20 {

              // group attributes:
              		:objectType = "gmi:LE_Source" ;
              		:gmd\:description = "Auxiliary LUT_CH4CIR algorithm lookup table" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "N/A" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2024-04-09T12:47:23Z" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "Auxiliary LUT_CH4CIR algorithm lookup table" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_OPER_LUT_CH4CIR_00000000T000000_99999999T999999_20151016T113037.nc" ;
                  } // group gmd\:alternateTitle\#1
                } // group gmd\:sourceCitation
              } // group gmd\:source\#20

            group: gmd\:source\#21 {

              // group attributes:
              		:objectType = "gmi:LE_Source" ;
              		:gmd\:description = "Auxiliary LUT_CH4RFC algorithm lookup table" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "N/A" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2024-04-09T12:47:23Z" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "Auxiliary LUT_CH4RFC algorithm lookup table" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_OPER_LUT_CH4RFC_00000000T000000_99999999T999999_20230720T134206.zip" ;
                  } // group gmd\:alternateTitle\#1
                } // group gmd\:sourceCitation
              } // group gmd\:source\#21

            group: gmd\:source\#22 {

              // group attributes:
              		:objectType = "gmi:LE_Source" ;
              		:gmd\:description = "Auxiliary REF_DEM___ reference data" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "N/A" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2024-04-09T12:47:23Z" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "Auxiliary REF_DEM___ reference data" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_OPER_REF_DEM____20190404T150000_99999999T999999_20190405T143622.nc" ;
                  } // group gmd\:alternateTitle\#1
                } // group gmd\:sourceCitation
              } // group gmd\:source\#22

            group: gmd\:source\#23 {

              // group attributes:
              		:objectType = "gmi:LE_Source" ;
              		:gmd\:description = "Auxiliary REF_SOLAR_ reference data" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "N/A" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2024-04-09T12:47:23Z" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "Auxiliary REF_SOLAR_ reference data" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_OPER_REF_SOLAR__00000000T000000_99999999T999999_20210107T132455.nc" ;
                  } // group gmd\:alternateTitle\#1
                } // group gmd\:sourceCitation
              } // group gmd\:source\#23

            group: gmd\:source\#24 {

              // group attributes:
              		:objectType = "gmi:LE_Source" ;
              		:gmd\:description = "Auxiliary REF_XS_CH4 reference data" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "N/A" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2024-04-09T12:47:23Z" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "Auxiliary REF_XS_CH4 reference data" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_OPER_REF_XS_CH4_00000000T000000_99999999T999999_20200710T082601.nc" ;
                  } // group gmd\:alternateTitle\#1
                } // group gmd\:sourceCitation
              } // group gmd\:source\#24
            } // group gmd\:processStep
          } // group gmd\:lineage

        group: subsystem_information {

          // group attributes:
          		:objectType = "subsystem_information" ;

          group: subsystem\#0 {

            // group attributes:
            		:Authors = "Tobias Borsdorff, Mari C. Martinez Velarte" ;
            		:Email = "T.Borsdorff@sron.nl, m.c.martinez.velarte@sron.nl" ;
            		:Institution = "SRON Netherlands institute for Space Research" ;
            		:Name = "Internal cloud mask" ;
            		:Reference = "To be written." ;
            		:Version = "2.6.0" ;
            		:VersionDate = "2023-07-20" ;
            } // group subsystem\#0

          group: subsystem\#1 {

            // group attributes:
            		:Authors = "Tobias Borsdorff, Mari C. Martinez Velarte" ;
            		:Email = "T.Borsdorff@sron.nl, m.c.martinez.velarte@sron.nl" ;
            		:Institution = "SRON Netherlands institute for Space Research" ;
            		:Name = "RemoTeC" ;
            		:Reference = "Hasekamp, O. et al., Algorithm Theoretical Baseline Document for Sentinel-5 Precursor methane retrieval, SRON-S5P-LEV2-RP-001, SRON Netherlands Institute for Space Research, 2022" ;
            		:Version = "2.6.0" ;
            		:VersionDate = "2023-07-25" ;
            } // group subsystem\#1

          group: subsystem\#2 {

            // group attributes:
            		:Authors = "J. Landgraf, O.P. Hasekamp" ;
            		:Email = "J.M.J.Aan.de.brugh@sron.nl, J.Landgraf@sron.nl" ;
            		:Institution = "SRON Netherlands Institute for Space Research" ;
            		:Name = "S-Lintran v1" ;
            		:Reference = "Landgraf et al., JGR, 106, D21, 27291-27305, doi:10.1029/2001JD000636, 2001" ;
            		:Version = "1.5" ;
            		:VersionDate = "2010-01-01" ;
            } // group subsystem\#2

          group: subsystem\#3 {

            // group attributes:
            		:Authors = "J.M.J. Aan de Brugh, J. Landgraf" ;
            		:Email = "J.M.J.Aan.de.brugh@sron.nl, J.Landgraf@sron.nl" ;
            		:Institution = "SRON Netherlands Institute for Space Research" ;
            		:Name = "S-Lintran v2" ;
            		:Reference = "Schepers et al., JQSRT, 149, 347-359, doi:10.1016/j.jqsrt.2014.08.019, 2014" ;
            		:Version = "2.3" ;
            		:VersionDate = "2015-02-11" ;
            } // group subsystem\#3
          } // group subsystem_information
        } // group variable_header
      } // group earth_explorer_header
    } // group ESA_METADATA
  } // group METADATA
}
